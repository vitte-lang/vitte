   d  x  �|                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �^Юn��P�P�Հ��P��p�P��P��c ��u�  �P��@K �        ^ݬݬݬ� � �!�社          ^�� �� ݬݬ�  �P[ЬP(@ݬ��-�  �P�@0Ь�@)ݏ�� ��'�  �P��P��P6��P�H   ���[P        ^��� #Џ,  �t� x�m� ~��N �P�b� #��U� x�N� ~��K� ��Q �P�=� ��7� ݏ�� ���           ^��� P��� P� �o������ P���� Ь@���       ^� ��� ݏ�� ��9�  ��w� P��o� ��Q� `��b� P��Z� ��@� `��M� P��E� ��/� `��8� P��0� ��� `���         ^��� ��
� ��� ���� ҬP�P��� P�P�� ��� ��ߗ ��ٗ ��� ��͗ ��Ǘ ��        ^ݬ�﹣  �P�ѼЬPѠ@� @  ݏυ ����  n��x� �� ݏ� ���  R��\� �Z ݏ�� ���  ЬPР<�<� � �m�  ��/� Q�P��P��Q3 ��� ݬ����           ^���� ��� P�PP�PP��� ݏ� �� �  E���� �� ݏ1� ���  )� ��  ��� �� Q�QQ�QQ�P�� �P���2       ^��� �Z ݏK� ��5�  Ï� �f� P�P�Y� ��W� PЏ�������G�   �   ^��0� P�PP�PP�PP��� P[�[W��� X�[X9�[Y�YX)�i��YW�i���giЭ�gЩ��Ч�Э���Y��WX�[W��[Z�Z��� !�j���j��ݭ�ݏa� ����  +�Z���U �[�� P�P~�[~��y�  �[�� �h  ^�ZЏ�����ڀ ��؀ ��ր �ͦ�XЏZ W�︀ V�ﳀ �變 P�@�s �J�{ � ݏ~� ��O "�J�{ ��x� P�@�s ݏ�� ���N �X�mP�XPݏ�� ���I  �P1��Zh�W}�� g2J�h Y�Y����1� ��� |� �)  �P�� ��� W��� ݏ�� ��tN @��� P�@��r ��� P�@��r ݏ�� ��GN �� ݏ�� ��2N �� �� �� Y	�Y��  J2I�^ Y2I�m P�P�u 1Џ�����h }�6� �9� ��+� P�YZ��U ��M 1��2J��o Y�Y�����1� ��( W� �(  �P� �� 2��	 ݏĆ ��~M ���~ P�@��q ݏ͆ ��aM ���~ ���~ Џ$d V2fP�P�����	2�P�PZ�V��V�f2fP�P�~ �2�Y�P1#�Y1�2�~ P1��J�y ݏՆ ��H  ��a~ P�@�iq ��Q~ P�@�Yq ݏ� ���G  U��4~  "��+~ �   ��~ ݏ� ��G  *��	~ ݏ�� ��G  ���} ݏ � ��G  ���} ���} �ͨ�P�XPn2hP2@�f P��   PY�Y(�Y��  2I��\ P�@�k � 2I�\ Z1��2hP2@��e Y��z} 2��~2h~ݏ� ���K �X�W��P1���P} 1� ݏ9� ���K ��<} P�@�Dp ��,} P�@�4p ݏR� ��K U��}  "��} �   ���| ݏV� ��pK *���| ݏ\� ��YK ���| ݏa� ��DK ��| 1U�Џ�����| 1o��P (�����I���| 1� �Yݏk� ��K �J�w ͜��ݜ�t��� �ݜ�P��� Q��� �Paݏ�� �ݜ�~��TB �ݜ�
6�͜�P��,��a� �	P��Z� Q��S� �Paݏ�� �	��B �͜��2I�h P�PP�PX�W[2I�h P�PP�PP�PP�PW�WP}`�� �Y͠�2I�g Y2I�f P2hQ�QP�Pͤ��ͤ���  �ͤ�P2@�Z Z2J�i P�YQ�PQ2I�Ef P2@�Z Z�͠�P1�� ���  � �;  1���YY ��WY 1���JY ��HY 1�� �v2  ��4Y ��2Y 1�Џa   ��1�Џa   ��1���Y �~�~�kݫ���V  �P��[2  1|���X ݏ{� ��+�  ��iO ���X Џa   ��� ��:  1F��X 1=��X Џa   ��1,��X Џa   ��1��X 1� ��  � ��A�  1�Џa   ��1�Џa   ��1��� �������P�� ��>X 1��k�� 1��� ��������P��� 1���X 1���kPݠЫ�Pݠ��T  �P͘�Ы�P�͘��Џa   � 1q�k��W 1g��kPݠЫ�Pݠ��MT  �P͘�Ы�P�͘��Џa   � 17�kPݠЫ�PݠЫ�Pݠ��T  �P͘�Ы�P�͘��Џa   P�P� �P��1�ݫ���?  �P�2� 1�� �k���<  �P�� ��OW �NW 1�� ݏ�������=  �P��� ��.W 1�� �k���=  �P��� ��W 1��k��n=  1�k� W ݫ���Z=  1kݫ���?  �P�� 1Wݫ��k��g<  �P�� 1A�kݏ������Z=  �P�s� ��V 1"ݫ��k��>=  �P�W� ��V 1��pV ��~V Џa   ��1���YV ��PV c���V ~���V ݏ�� ݏ\2	 ��*I ��(V �ݏ\2	 ��& �P� ��������P�k��S  �P��d/  ݏ�� ����  ���U Џa   � 1j���U �kݫ���xS  �P��+/  ���U ��U 1AЫ��� 16��U �kݫ���DS  �P���.  ��U �U 1��U ݏ�� ��;�  �k	�k�@   ݏ· ��!�  �kɏ@   k~ݫ�ݫ����R  �P��.  ���� 1���,U ݏ� ����  ݫ�ݏ�����kݏ�c ��1O  ���� 1|��� 1s� �k�������P�� 1\� ݫ�ݏH   ������P�� 1@� ݫ��6������P�s� 1(ի�ݏ�� ���  ݫ�ݫ��6��W����P�H� 1��k� ���@����P�1� 1�Ы��&� 1�1e�1y���Ы��� 1���� ݏ� ����  1���T ݏ/� ����  � ݫ�� ��������PݏH   �������P�� ���S 1j��P� ݏS� ���  1R� ݫ�� �������PݏH   ������P�t� ��S 1#��S ���P��c ���PЏ@   �c 1��k��??  ��pS 1��k��,?  ��]S 1�Ы��� 1���5S �kݫ����P  �Pk�P��,  �kPݠ@���A  1��kݫ���P  �P��O  1����R ��S  �P�kݫ���P  �P��=,  1^�k��iG  � ��E  1K� ��E  1A�k��LG  15� �K  1+� �J  1!��R ���V  ��R ��|R ��sR ���V  ��fR ��� ��� ��� ��� ��ۈ �JR 1���9R � �G5  � �tV  �ﶈ ��� ݏk� ��^�  � P� ��R `� P��� ��a� `1mݫ��ﷃ  1`� �+  1Vݫ���|$ ��MH 1Bѫ������ݫ���^$ ��/H 1$1!� ������H ݏ|� ��y�  ��H � �/�  �P��� � �!�  �P��� � P1Vݏ�� �  ��� ���# ѻ�Ы�Pՠ<��� ݫ���z�  1Ы�PЫ�D��}� ��6o  �Pݫ�ݏm   ��LX  �P�ￂ  1� ѻ�)Ы�Pՠ< ��J� ݫ���$�  ��6� ��k# $��'� ����  � �]�  �P�f� �P��E# 1� ѻ�4Ы�Pՠ<+���� ݫ���ο  ���� �/� ��)� ��
# Tݫ����  �P͜���� ��ln  �Pݫ�ݏm   ��W  �P����  �͜���� �́  �P��� �P��" �P ���l�1��1r��0� P1� ݏ�� ���  ��I� ���  1� ��<� ��0� ���  J��4F ��� ��O" ݫ����m  �P� ݫ�ݏL   ���V  �Pݏm   ���V  �P��=�  z���� ���� �  S���� ���E ��� ���! ݫ���Xm  �P� ݫ�ݏL   ��lV  �Pݏm   ��]V  �P��Ѐ  �P �+���1���^� 	��U� 	��\E ��TE ��6� ��o! � �����13��!� ��V! ��� ��E Ы�PЫ�Dݫ���l  �P� ݫ�ݏL   ���U  �Pݏm   ��U  �P��+�  ���� ���  ���D � �����1�1�ի�Ы�PЫԠDݫ����  ��D ݏш ����  � ������ �  �P�d� � �  �P�R� ��cD ��� P1zݏ� ���  � �u  �P�~� �P��]  ի�	��� [ѻ�Ы�Pՠ<��� ݫ���ۼ  ԫ�6ի�	Ы�PЫԠD���� ��k  �Pݫ�ݏm   ��T  �P��  1� ի�	��� 9ѻ�Ы�Pՠ<��� ݫ���o�  ԫ�� �~  �P���P��F�  � �~  �P�� �P�� 1� ի�	��L� bѻ�Ы�Pՠ<��4� ݫ����  ԫ�=ݫ���?�  �P͜���� ���j  �Pݫ�ݏm   ���S  �P��J~  �͜���� �!~  �P�*� �P��	 �P ���s�1y�1���� ��� ��� ��B ի�Ы�P��� �Dݫ����}  ��Q� Pqݏ� ��=�  ݫ���;�  dի�
ݫ��� ի�8ݫ����i  �P� ݫ�ݏL   ��S  �Pݏm   ��S  �P��w}  
ݫ����  �P ����������� ��, ���� 	���� 	���A ���A � �����1����A ��� �  ݫ���� � �e������ ��� ��� 	��� ��A ���b���1w��a� �����ݏ#� �  $��]A Ы��C� � �l�  ��.� ���  ��(� ��� m��(A 1��� �����ݏ1� ��G�  Ы���� � ��  ���� �ﱐ  ���� #��MJ Ы���� � ��  ��Ā �  ��@ ݏB� ���  ��@ 1�
��� �� � � ���[Q  �P͜��͜�P�͜�Q��R�R�͜�Qˏ�����S�SR��͜�PѠ�P   ��B� P��c ݏX� ��r�  Џv   ݜ��͜�Pݠ�͜�Pݠ�͜�Pݠݫ���kq  �P���͜�Pݠ��LP  �P͘��͜�P�͘��ݫ��͜��:��P  �P͜��͜�PЫ��D�͜���
{  ��'I �� ��n�  ��? 1�	�� ݏd   � � ݏa   ��rr  �P͜��͜�PЫ��l� ��f� �@��͜���3"  ��P� P��=� �c Ы��4� � �]�  ��.� P��c ���  1d��� ݏd   � � ݏa   ���q  �P͜��͜�PЫ��@��͜����!  ���> 1�ݫ���������> 1����> � ������� 1�� ������> ݏ}� ���  � ��y  �P�v� � �y  �P�l� � �y  �Pﲿ �P�� ��b> 1WЫ�PЫ�D� �y  �P �P���e  �Pݫ�ݏm   ���N  �P��py  ��> 1��> � �;y  �P�D� �P�ￍ  Џ�����.� ݫ��� ���= 1�� �3����� �� � ݏw   ��p  �P͜�ݫ��͜��:��wN  �P͜�� ��x  �P�|� �͜�PЫ�D�͜����x  � �x  �Pﱾ �P��,�  � �������[= 1P���F  ��F ��F �F 11�k��Xp  �P�i� Ы��F 1��X� 1B��qh $��hh ��_h ��Vh 	��Mh ���| ݏ�� ��=�  �kݫ�ݫ���M  �P��� 1��;������h ����h �����g 	���g ���1h����g 	���g 1S�����g 	��g 1<�1{���g 	��g 1$�1c�1`�1]��kݫ����~���L  �P�V� 1��������kݫ�����L  �Pݫ����L  �P�"� 1�ݏ ��>�  1��1�����kc  �Pݫ��k��L  �P�� 1�� �k���~��kL  �P�Լ 1��kPˏ�����Q�Q�@   �kPˏ�����Q�Q�`   ݏ� ��Ʋ  �k �1D�� �kݫ���L  �P�u� 1*����b  �P�kѫ��N   �~�	~���K  �P�E� 1��k��	s  �P�2� 1��kݫ�ݏr   ��K  �P�� ��� PЏa   �<Џa   ��� ���� PР@�� 1�ݫ���r  �P�ٻ 1�ݫ�ݫ��6��WK  �P��� 1uݫ�ݫ�ݫ���K  �P僚 1[� ݫ�ݏH   ��!K  �P 1?ݫ�ݫ�ݏF   ��K  �P�m� 1"ѫ��D   -ݫ���a  �Pݏ� ��q�  � ݫ�����J  �P���k��� � � ���J  �Pݫ�ݏE   ��J  �P�� 1��k�� ��"C b��� P��c Q��� P��c ݏ0� ����  �� �� � ݏa   ��]l  �P͜��͜�P��Y� �@��͜���&  � � ���J  �P�~� �kP�� � �c 1$� ���`  �P�\� ��V� P��� �<��G� PЏ @  �@�k(����B  �P͘���&� P�͘����� P�͘��1�� � ���I  �P��� ���� Pp�� �1�� ��3  �P�۹ 1�Ы��й 1��kݫ���?  �Pﺹ ���� Џa   ��1`ݏ����� �������P 1E� ݏ����� �������PݏH   ��s����P�d� 1� ݫ�ݏH   ��W����P�H� 1�1��1��1��Ы��4� 1����P��c 7�� ݏD   � � ݏa   ��j  �P͜��͜�PЫ��@��͜���  Ы��� � � ���gH  �P�и ��� P��n� �c 1r�P��   j�{���������$�-�>�O�jY�l�w�jj���j��������j�3�jjo�����jj�������)�H�jjd�{� �)�4�j]�������*�B�m��������� ��G�n��jj��j��j������jjj)�5�jjjj?�I����
�j�(�F�I���7��������M�������jjjjM��������X����9�jT�j]�_������������������&�>�A�D�_�a�c�e�g�i�k�m�����j������&�(�@�p����������+�H���F���������
�%�Q�m�p�s�v���1��     ^Ь[ӏ@   [$ˏ����[~ݏh� ݏh2	 ��72 Џh2	 P
�K��u P        ^ԭ�����[x�����[խ���[PxP�� �[�[�1��K�Z�j-1O�Z�j�X��Z�j1;��� �jP1� ��� 1#��{� 1��v� 1��� 1���{ 1� ��u 1� ��2� 1� ��5� 1� � 1� ���t 1� �ﲊ 1� ��)� 1� ���u ��
� 1� ��я ���� 1� ��u 1� ��u 1� �j~ݏ�� ��j�  }�P�B   8\�������������������������e�I�������������R�������������������������n���������w�����������������������������������1q�1��1� �K�P�`-1� Э�P֭�{� ��Z% � �K����- �Pi�K�ݏ�� ݏ�� ��T' ���7% ݏ�� ݏ�� �K���' �P,�K�ݏ�� ݏ�� ��' ����$ 
�P ������[1�����t( �P��� ݬݬ���  �[�[�p  �[P��c �[�� �  � ��  � ��  � �������z� ��t� PԠ@��j� P����_� P� ���T� P� ���I� PЏ@   ���:� P� ���/� P����$� P��0��� P��4��� P� �8��� P� �<���� ��2 � ����� ��'  � �#�  ��}� �P�P       ^��Us 1� ��	 �Is �[�
��?s ��\! �PZ��0s Z�[+�Z�j�	 �j��s ���   ��	s P��s �`P1� ���r ��r [�[���r ݏt2	 ��3+ �P��r �[�   ~��t2	 [��r ��r � ���, �P[Џt2	 �r ���r Џ����Pk�[�r ���r 1;�ݏ   ݏt2	 � ��, �P[Џt2	 �]r ��Wr Џ����P'Џt2	 �Cr ��=r [P�`��3r P��,r �`P        ^Ь[��� P�P�P�� Pݏ� ���� ݏ� ݏН �� �kP��� �[�k�[ݏ� ݏ� ���       ^Ь[��Z��Y�YP�Z@��� �        ^Ь[ЬZ��� Y�[i��oq ��gq P��`q �`P� ������P[�[P�Z@�� �Y�7 �Y�[i���-q �Y�Y� ��S�        ^�ݏ� ��L����ݏ"� ��=����ݏ-� ��.����ݏD� ������ݏK� ������ �s� � �&  �Z�Z��   Џ� J��� �Z�Џ� [2kP�P�[@��� �k�[�ЏT� Y�i��P�PЏ� @��� �Џ�� Y�i��P�PЏ� @�� �Џ�� Y�i��P�PЏ$� @�� ���� � �|          ^Ь[�X���o ���o P���o �`P� �|����PZ�Z�:� 1��ZP1�ݏ�� ���  1�ݏ�� ���  ��� 1����o ��o P��o �`P� � ����PZ�ZP1� ��y� 1q��ZY1��
Y1��Y1��Y1��	Y1��Y1��Y1��0ZY��Bo ��:o P��3o �`P� �����PZ�ZP�@�l� `�YYP�PP�PP�0ZQ�QPY���n ���n P���n �`P� �{����PZ�ZP�@�(� �YYP�PP�PP�0ZQ�QPY��n ��n 1� �P
�l   &�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�Y�Y�Y�Y�Y�Y�Y�Y�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�/�A�/�/�/�M�/�/�/�/�/�/�/�5�/�/�/�;�/�G�/�S�1R��ZY�YY��� '8��Y��Fd  �PY�X	�Y�� x�� �� ˏ ���YP�P�� ;��;� (�[�X[�Y���(  �X[ݏӞ ��ӣ  �X�Y��	 �X1<��P�����1f��P
1n��P�\   1x�1V� ��v� "J���� �[�X[	� ��}(  ,�X~�X� ��]	 �Xݏ������N	 ��8� P�X@�+� 8�Xݏ�� ���  �X��k ��k �Xݏ� ���       ^���l ��yl P��rl �`P� ������P[�[PJݏB� �  S��I� H��Al ��9l P��2l �`P� �����P[�[/ ��l �P�������P
��P*��1u�   �    ^���k ���k P���k �`P� �f����P[�[P�@�� Z2�P1���k �[��k 2��� ��� �� 2�P1��[ݏY� ��Ҡ  1�Џ8 �� ��[������� ��  �P[��W�  �[P1��[1���3k ��s� ���3 	Џ@   ~��3 �~�~ݏ8 ��X �P�� �PW�WP���c PY��=��t3 5��h3 �g3 2�~2�~ݩ�������P�
� ��� �� �!P1��63 	��*3 P�P�P�"3 �W�ת ��� �Ъ �P1���� Џ8 �� ��[��������Xj ��Pj P��Ij �`P� ������P[�[P1q��b� 0��Z� ݏy� ��f�  ��[��{���Џ: X�hWx�	� �� �hP��� �hP�0P�P��� ,�hP��� �hP�7P�P��� �hPW   P�P�� �X�ӏ  ���� 	��� ��٩ 1j��[��������yi ��qi P��ji �`P� ������P[�[�e   	�[�E   b��Ci ��;i P��4i �`P� ������P[�[+�[-��I� P��B� ��e`��i �[��h Џe   [��[��Y������h �[��h ��h ݏ8 ��^ pP��� ��� �� �P1��h �[��h ���� 0+Џ9 X�hx�� �� �hP�0P�P�� �X�1��Џ8 X�h�
�k� P�hQ�QP�0P�\� �X�ˏ�  �M� V�V	�V� �����u� ��l� ��h ��h P��h �`P� �����P[�[�L   	�[�l   	��/� ���g �[��g ���� �� �P1+�P.11��P�E   1f��P�X   1o��P�e   1N��P�x   1W�1�����g ��zg P��sg �`P� ������P[�[P�@�� &��Pg �[�Ig Џ8 �r� ��.�����1����/ 1n��"�� ��� �d� �P1v�'�g� ��� � ��������>� ��� �7� �P1I���f ���f P���f �`P� �X����P[�[*1��� ����1�勵 � �  1 ���f ��f P��f �`P� �����P[�[=1��ЏQ   ﰦ ��^� 辶 �P1���Mf ��Ef P��>f �`P� ������P[�[-ЏO   �k� ��� �d� �P1v�[>1N���. ЏE   �@� ��� �9� � P1K���e ���e P���e �`P� �Z����P[�[+1��ЏN   ��� �料 �� �P1���e ��e P��e �`P� �����P[�[&1����i� ﴥ �贈 � P1���Me ��Ee P��>e �`P� ������P[�[�|   1k���� �h� ��]� ��W� P1o��e ���d P���d �`P� �~����P[�[<Џ@   �� ��ͽ �� �P1*�[=1�ЏR   ��� �墳 ��� �P1���d ��d P��d �`P� �����P[�[>ЏB   ﶤ ��d� ﯤ �P1� �[=1��ЏT    ��@�  �P1� ��/d ��'d P�� d �`P� �����P[�[PЏP   �M� ���� �F� �PY16��P=���[ݏ�� �神  .�P A�S�X�'���������J������7���4���7��$�'��ݏ�� ��k�  1��       ^Џ� [�kZ&�jPʏ����P��h ��Pʏ����P��� �[��Y�Y���Y���Y *��h ֭���h �� ֭쐭�� �Y�Џ� [�kZ9�jPʏ����P��h PxPQ�QP��Qʏ����Q�� Q�QP�� �P��[��YЏ � [�k*����ޭ�P(k`�[P(`kޭ�P�[Q(`a�Y�[��Y����Џ� [�kZ2�Y�� ���� �[֭��        ^��� 
Џ����P1���� Pʏ����P��h P�PP�PP�PP�PP��d� Qʏ����Q�� Q�QPˏ ���P[	�� [
Џ����P1_�[P��� PZ�jݏ8 �� �P1%2�P1
��\* �[* 2�~� 2�~�������P��� ������a �!P1�2��ޡ ��ء P1�2��̡ �"P1���* �︡ �#P1����) �嵐 �#P1����) �1 � P1���#a Џ8 �\� �� �������a ��a P��a �`P� �����P(1Џ8 �� �� ��N������` ���` P���` �`P� �U����P"1� Џh ��� ���` ��` P��` �`P� �!����P[�["C�[
	�[�����1� ��� P��� �[`��� �/ ݏ�   ݏɟ �  �Џ8 �g� �� �������"` ��` P��` �`P� �����P)��&� P��� �`�;PLݏ؟ ��/�  �P;ݏ� �  �P ��.�@�N�b�v�����Z2�P�P[1��Џ����P         ^���_ ��_ P��~_ �`P� �
����P[�[#�[�������[_ 1Џ8 �� �� ������Z��:_ ��2_ P��+_ �`P� �����P[��� 1�
ZP�[P�0PZ��_ ���^ P���^ �`P� �����P[����^ �Z�Է Џ8 ��� �� ��.������^ ��^ P��^ �`P� �5����P[�[
IЏ� Y�[����^ ��}^ P��v^ �`P� �����P[�[
�[�Ҕi�[�������L^          ^� �l�  ݏ� ݏh ݏ� ݏ�� ��A�  �   ^Ь[�[1�[� 	�[��� ݏ� �ﵓ  Ы@��խ�ݏ� �  ���P���c PZ��c Aݭ��jݏ�� �� ݫ��QV  ��& ݫݫݬ������Pݏ� ��t ݬ�[��%  ЫY�Yݬ���&  �P�ЪX��	����c jݏ � ��6 �Y���U  ݬ��7����Pݏ.� �� ݏ4� �� �X��U  ݭ�2�~2�~��~�������PݏF� ��� �X�@   ��1W�X�XJ��<% >�X9ЬPӏ@   ��jݏa� ���  �P�������������������1�YX1�2�VЫ���Y��ӏ`   ��oˏ������P�P�`   D�F��� Э�P�@��� F��� #Э�P�@��� Э�P�F�s� @�m� 1c�V֭����P�Pˏ������Q�QP���ѭ�ѭ�	ѭ�
2�P�P�Ѭ
Ѭ	Ѭ1��W��a �W������Pݏ�� �� ӏ@   �*� �ˏ�����~�Z��-  �Pݭ���  1x1�ЬP1��WPխ�1a)1\�P����" ��" " " " " " " " ��" " ����1z�W�W(��#  ��ˏ����YP�P�@   Э���� 11E�W�W1�15�W��ݪ���  1�1�W�1�1�W�W1�1 �W ��ˏ����YP�P�@   Э� 1�1� �W�/ݏ�c �Z��0  �P1� Ѭ���" ݭ���  1\1� �W� ���" P���" ѪP1� ݭ���w  x�W ��ˏ����YP�P�@   Э��� 1Q�W�I2�P�@�C� 1�7�W�W1�(�P��o�����������L�����L����$��������ѬѬӏ@   �1� � �
��y� P�PP�PP��0� P��ս�k���P��c 
]���P��c O���P� �c ;���P�j�c +���P2�c ��խ�έ��ݭ��jݏ�� ��Y�  ����߭����$  �PZ}��l! ��>Ѭ8Ѭ2Ѭ,Ѭѭ� �Z���&  �P���P�@���P���c PZ52�~�jݏ�� ���  Ѭˏ����YP�P�@   Э� 1���?^ ݏޡ ��\ �Y�jݏ� �  �Y����ѬѬ�P��  P�P�	Џ'������� �Ѭ
ѬѬ3��c� �� ��0���ݏ������#���������ݭ������)ˏ����YP����YP����P��P������谫�ӏ@   �#� � ˏ�����~�Z��<  ݭ����  1� ЬP1� ݏ � �Z��)  1� � �Q  �P�ˏ����YP�P�@   Э��B� 1� � �tQ  �P�Ѭ� ��iP  ݪ��O�  1� � �MQ  �P�~ݏ�c �Z��  Ѭ��| ݭ���6  W��j ���b ݭ���  =��t� ���4 ��
&�P7���I���I�p�p���" " ��" " ��" ������� �d   ݏd   ��� ݏ � ��/�  ��	��Э�P�@�� �Э�P�Z@�� ЬP��	)��	$�P��      ����            ��    �����[ ݪ2�~2�~ݏ!� ���          ^���� 2�2��� ݏF� �  ��׹ P��й Ь@�Ϲ         ^� ��  ݏ�  ��~� ݏb� ��I�  ��k� P��d� Ь@         ^��aT ������ �i  � �t�  �� � ﯌  �� Џ�����.T ��(T �� ��� �� ��� ��� ��� ���n D���S �p� ݏ�� �金  ��ƭ ݏ�� �  ���� ݏ�� ��z�  Џp� �S � � ��x �� � Џ�  ���M     �   ^� �� ��"Z ݏ�� ��> �[�[�U� 1� �K�Q� Z1� �ZP���c PY���Y (�Z�iݏ�� ��� ݩ��L  ݏɢ ��� ѩ)�� �� � ݏa   ���E  �PX�Z�@�	�X�������=Щ��Џ'�����	�ݏ�  �Y��]  ЩK�� ЩK�o� ��Э��!ݏ�  �Y��1  ЩKﴶ ЩK�C� �[1���H� � ��L  � ��>�  ��T� ��5� P���c PY��	��ݩ��J�  	�Y���h  ЩW�WP�Pˏ����WQ�QPW�W�W	�P�P�P�� ��� 2�~2�~��DP  �P��ͫ �i��Ŷ ݏ(� ��g  � �)   �﫫 2�~2�~�W��  �P[�[��h         ^�[�[�v� |�K�t� P���c PX��`�K�^� �A� � � ���"  �PZШ���K�m� ��	�� � ����!  �PY�Y�Z�:���!  �PZ�Z��JL  Э�����[1{�        ^Ь[ЬZ�[P���c PYЩPv� � � � � ݏa   ��C  �PX�[�@�Z�P�Z�	P�
P�P��Z�
~�Z�~�~�X��D���3�Z,��Z#��Z��P	������      ���� � 2�~� ݩ��D���       ^Ь[� � �� � ݏa   ���B  �PZ�[�@�[��Z�����     ^Ь[ЬZ�[1� �/ݏ� ����  �P��Џ� �����ݭ�ݏ�B	 ��� �"ݏ�B	 ���  �P��������� ���� ��X� ݏ�B	 ݏˢ ݏ�B	 �� ݏ@   ݏ�B	 ��|�  �P���  �P[�� ��k����� ��^����� ��Q����� �Z�x � � � � � ݏa   ���A  �PY�[�@��T ��: ���
�Y�����7��3 �� �	���Y��v����� �
���Y��^���Щ@[�[�������[�[P��[� �c ��G� P    �   ^Ь[�[P�@�\� Y7� ��� ��X���ݏ������K������B����� � ~��4����YP2�c ����T (ݭ��Y�YP��c ~Џ� ~ݏԢ �� ��? �P��1 �	P�
P�P���KＧ � �� � �[P�@ �� ���P��Ɏ @��� �Xԭ�Э���[Y�Y�A� 1� �I�i� V�V��o����V	�V�p  ݏ� ���  �VP���c PZѭ�
Ѫ��Ъ��Ѫ��Ъ����z2�~ݪ��  �PW��@���Pˏ����P��2�~2�~ݪ��;  �P��խ��jݏ� ���  ѭ��# Э�� �WXP�WP�PXP
�WXP�P�WPX�Y1�ݏ��������X�� P�XP�P�� P�X�� P�P�XP�� ѭ�
=���ݭ�� ݭ���  �P� ݭ�ݭ����  �P��Э�X���PЭ�@�R� �� ݏ(� ��-�  Э�P��g @�-� ���P�X@� � ���P�[Q�A�ܥ @�
� ��tR 1� ���P�@�� ���P�@�� ���P�@�ڌ Э�P�@�ό ���~���~���~ݭ�ݏ=� �	�L ���P�@��� Y�I��� '�I��� �I��� P��c ݏa� �� �Y��[P�@�4� � �[��� ݭ�� ݭ���%���         ^ݬ ݬݬݬݬݬݬݬ���           ^� �L���        ^Ь[�[P���c PZЪP-E�jݏq� ��Ȁ  �Z��  �P[�[P���c PZ�P ��P��P��P�@   �����	��[��I���     ^Ь[ЬZ�Y�YI�Y Q�YQ[Pʏ����Pݏ�� ��ɀ  � P}�P ��P ��P�@   ��P�`   ��Y�ˏ����[P,�ZP�@�� P@�P;� P6� P1� P,�P'� P"�P�����������������������������       ^Ь[�Y�Z�ZZ�Z Q�ZQ[Pʏ����P'ݏ�� ��  xYP1� ЬP֬�@��� Y�P ��P ��P�@   ��P�`   ��Z��[
� PC�[ݏܣ ��7  ЬP�@�<� ݏ� ��  � PЬP�Y@�� Q�QP       ^Ь[��]� [1� ��Q� [�[��F� ݏ�� ���~  �[�2� 1� ��)� Z� ZP� P�PZP
� ZP�PxPZ�Z[��� [Y�Y��\  M��� ZY�Y���[  ��� [P� PY�Y��[  ��ͮ [Y�Y���[  �Ｎ [ݏ� ���~          ^� [Ǭ[PĬP�P[PǬ[P�PŬP[�[�����        ^��G ݬݏ&� �� ��P���c P[���ul ��� 	��� ��\l ��Vl Pn1� 1� ˏ�����P�P�`   �P�P�P�N ��N ��sA  2�~ݫ�������P���  ��	��ݫ��6�  	�[���]  �P����������      ��� ��M ���� ��u� 2�~2�~ݫݬ��           ^ЬZЬ[��F �[ݬݬ�Zݬݏ=� ��i  ��s� Џ� �f� �$�]� ��W� PԠ��M� PЬ���A� P�Z���6� PЬ���*� PЬ���� PԠ��� P�Z��Q�A�V� Q�Q�Q����� P�[� ˏ����ZP�P�`   ,ݬ��~�ZP�Pˏ����ZQ�QP~��:����P��� 1��P��@�c ��P��c Pʏ����P�P��� ���� ��fj 	��]j #ˏ����ZP�P�`   �ZݏW� ��{  ˏ����ZP�P�`   �ZP�Pˏ����ZQ�QPZ֬V�ZO��� PРQ�A�^� ���P���c PY����@�ݏ}� ��{  ЩZ2��2����[1-�        ^��i ��i 1� ��� PѠ��� PѠ���� �� s��y� Pˏ������Q�Q�`   Z��� � �  ��R� Pݠ ������$�@� P�P�� ��0� PР�Q�A�x� ~�~������� ��  �P1� ���h 	� �������i �~�~��$>  �PZ� �?  �P[�[����  ��|� � �������- 	��}J ~�Z~���=  � � ���o  �PY�[�@�YP        ^ݬ��%+  �P[��[��CW  �[��:|  � �s    �    ^��9C ��� ݏ�� �� �  ��h P	��h 11�P���� ��Џ� �� ��� PР[���� PРZ���� PРY���� PРXˏ����[P�P�`   t�J�� W���� ��������� �Z� X�WX�Y�Z�[������P�������WX�W�WX�W�Xݏ�� ��x  �XݏϤ ���y  �XJ��� N�[�[	�Y�Z�[������P��v���,�X�Xݏ� ��dx  �Y�Z�[������P��H������ � ������ ���f �    ^Ь[���\ 1���f 1���f 	��f ݏ� ���w  Џ�����f 1���f 	��yf ?� �N  ��}� PР�t� �[� � ���=  �P�:��2  �P[�[��<  1f�[1_��H ݏ&� ��sw  1>��A �[ݏ1� ���  ��� PРW��� PРY���� PРX��� 	��� Z�X�Y�W��U����PZ��̿ Pݠ ������[�X�Y�W� � ���3  �P�:��y  �P[Џa   �<Ы@�<ԫ@ݫ<��L  �P�<ѻ<Џa   �<Ы<PР<�<Џq   k�[��mL  �P[ѻ<�ZЫ<Pp�~��T  Hѻ<ݏ=� ��nv  �Z�Ӧ ,�Z �Zݫ<���S  �[��L  �P���;  �Z復 � �
   �[���x  �   ^��վ �� 1%��ž Pՠ��F �$ﲾ �מּ PР[�[M� ��ֽ�н�Z�J�߀ X1� �XP���c PW��s� P�� �~2�~2�~ݧ�X�����1� ˏ����[P�P�`   1� ��:� ��ֽ�н�Y��+� PРQ�YA�r� ��� �� d��� V�� � P�VYQ�Q� ~��� Pݠ��� P��~��ڽ P��Q�Q��ʽ Pˏ�����R�RQ~�ﶽ Pݠ������1��      ^� Z� �� `� PР[�[ˏ����[P�P�`   4��^� Pՠ��R� Pՠݏ\� ��t  ��7� P��	�$�)� ��Z� �          ^��> ��� ݏf� ����  ��D ��D 7��� �� *��ռ Pՠ��Ǽ PԠ� �����	�$ﳼ �     ^Ь[ЬZ�jY�[YP�[P�PYP
�[YP�P�[PY�Y襁 P�P�%��� ݏ�� ��%t  ݏ�� ��t  ��Yj�YP    �   ^Ь[ЬZ2�~ݫ�������PY�jX�X��2�~2�~ݫ������PW��@�X�%� P�PWݏȥ ��s  �WX���Y��P�YP�P��P�Y��P�P�YP��έ�XA��	*� WP� P�PWP�WP� PW߭�� xW~�������PX߭��Y�W�������PX��ѫ�'����X��X��PЭ�j�P  �    ^Ь[ЬZլЪPЫP�PWլЪPЫPRլЪP2�P�PV�VP�@�W} Y�F�O} XJ�Y�XB�Y�X:� Y� X2ݏ� ��r  � Y �P���������������������������ѬX�Xݬݏ�� ���q  �X�լ>�Y� P�YP�P� P�Y�� P�P�YP�� լݏ� ��q  �P1� �Y�� P�YP�P�� P��P�PX'�Y� P�YP�P� P�Y� P�P�YP� լ+�� �(� P�P�ݏ� ��q  ���h �P^Ѭ!ѫ�V ��Pɏ@   �Q�PQ�P7��7 ���/ �γ P�P�ݏ4� ��Rq  ��� �W��P       ^Ь[�Y��� Z8��� �Z*��� ��� ݏO� ���p  �Z�Z�Y�Z�[�������Z�Z�Y�Y
ݫ@��VQ   �   ^Ь[ЬZЬY�[���Z���Y���V�X�Wԭ�ѭ�1� ޭ�P����Q�QQ�QP�`PYݏ[� ���o  �P1� j�V��V^�W�ޭ�P����Q�QQ�QP�`WB�X�ޭ�P����Q�QQ�QP�`X&�P���������������������������������֭�1]��X�X.�X�V�W1_��W�P�P%�X�W1C��W�WX�V�
XP�XP         ^Ь[ЬZ�k!ݏt� ��o  �Z�P1� ��r? 	�Z��1  Ы����y ��Z��   Ы�ЫYЫXӏ`   Y:ˏ����YP�P�`   �XP�X�@��y ����YP�Pˏ����YQ�QPY�ݪ��:  �P�ˏ�����Y�Y�Y		�Y
�Y��ZP      ^Ь[�kZЏa   k�Zw��P�PP�PP� Pˏ�����Q�QPX�Z�H   � X�Z6��@   XЫ@PР<YЏa   �@Ы<P�X�ݫ<������Z6	�Y�﹞��Ы<PР@�@Ы<PР�  �    ^Ь[ЬZЫX�X1^ˏ����XV1� �XP�Pˏ����XQ�QPY�VWˏ����YVc�W�`   �V�@   ݏ�� ��Nm  �X*�W�@   !�V�`   	�V�@   ݏ�� ��"m  �X�YP�Pˏ����YQ�QPY��Z��0  ��2  �	Z�Z	�Zg��  ^�X�XTˏ����XP�P�`   ֫������X7ˏ����XP�P�@   &ݏĦ ���m  �XP�PP�PP� Pˏ����XQ�QPX��� 7ˏ����XP�P�@   &ݏ� ��Zl  �XP�PP�PP� Pˏ����XQ�QPX�X�     ^Ь[ˏ����[Z�Z
�[P�P[�Z�[P�P[�[P       ^Ь[�[�P�[�P�[�P�[P      ^ЬZЬ[�Z:���� �Z,���� �Z���� �Z���� �	Z�Z��� �Z�Zݏ� ��ek  ˏ����[P�P�@   A�ZPݏ>� ��Bk  �Z*�P�������������������������������������ӏ@   Z��?� ݏa� ���j  �ZP1��ZP1Q��� ݏx� ���j  �ZP1_��� ݏ�� ��j  �ZP1C���� ݏ�� ��j  �ZP1'��� ݏ�� ��j  �[���B  �P�ZP1� ��� �	P1� �P1� ��� ݏƧ ��?j  �ZP1� ��c� ݏܧ ��#j  �ZP1� ˏ����[P�P�@   ݏ� ���i  P�[P�Pˏ����[Q�QP[ˏ����[P�P�@   ˏ����[P�P�`   ˏ����[P�P ݏ� ��i  �ZP;�Zݏ5� ��j  *�P>���������>�>���Z���������v�����v����     ^Ь[�kZ�ZP���c PYթ-�Z�Z�p  �ZЏ�c Y�Y�ZkݏG� ��i  ΐ!�
�kP��c i�Zk��9 �Z�k�iݏY� ���  �YP         ^Ь[��
Pˏ����P~�k����  �P���c PZѪԪ�ZP&�Z[ժ�Z�Z��� Џ�c Z��ZP         ^��� � ��`        ^� �$a  ��� P�@�ʘ [�[�[��a  Ы[�� �sa  Ѭ� ��`  �ZЬP�@ [�[1� ��8 #��	~��
~Ï�c [P�P~�kݏ�� ���  ѫ��Ѭ�kݏ�� ���g  ��
	�[��>  �[�������PY�Y[(ki��	PѬP�[YЫ[�Z��YZԫЫ[1e�ЬP�@�� �ZE��
~�j���  �P���c PY�YZ(jiԪЪZ��P�@ﶗ ���P�Y@輪 �     ^Ь[�[Z�Z��� Џ�c Z�Z[ݏ�� ��ug  ժ�Z�(kj��
����
P�P�
��0 �kݏ˨ ���g  ��97 %Ï�c ZP�P~Ï�c [P�P~ݏ� ��>�  Ï�c ZP�P�>� ��8� P      ^Ь[��
Pˏ����PY�[Z�Z��c 	Џ�� Z�Z�Z[J��
Pʏ����P�PY8�kj3��
��6 %Ï�c [P�P~Ï�c ZP�P~ݏ�� ���  �ݏ� ��if       ^Ь[�[P
�P&�P!�P����        �����[P        ^Ь[ЬZЬYݏ�� ��e  �Y��h  �Z�[�6��     �(   ^ЬYЬ[ЬZ��)> 4Ï ZPǏH   P~Ï [PǏH   P~�I��S ݏ�� ����  �Y6� �Z�[�������P������1lˏ����I�U ���Y�L   �k��. ݏʩ ���e  1Z�Y
�kr���[P1#�YD�k?ѫ@� @  5Џa   kЏa   jի<ݪ@��g  Ъ<P1�
ݪ<��g  Ъ@P1�
�Y�Y�k�jѭ�1� �k��j��YP���- ݏ� ��Te  1� �P�V   ����� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��������������������� � � � � � � � � � � � � � � � � � � ���Y�m   �Y2ˏ�����Pˏ�����P�P ݏ� ��7c  
�P��������Ն ���[իDѫD��ЫD���ZժDѪD��ЪD���� ��Z�[�Y��  �PX�X��   �P��ӏ@   ��ݨ<��  �Pݏ� ��b  ӏ   ��ݨ<��)  �P�<B���<Э�P(ݨ@��  �P�@ӏ@   ��ݨ<���  �P�<�P��
 
 
 ������Y�r   ���+ 	�X��	  ���"���Ш<PШ@P�PWЧ�Ч�Ч�ӏ   ��ݏ   �X��p  �PXӏ   ��ݏ   �X��T  �PX� ���X���  �PXӏ   ���X��d  �PXӏ @  ���X���9  �PXӏ   ��1�Ш<[Ш@Z�YP1���1� P���c PVѦ7�fݏB� ��Wa  �P�P��P��P����� �@Ԩ<� �X������1\Ц�2��2��ѨЏ @  �@Ц�<Ԩ�
��hy��P[Џt   hЏ @  �@���<\Џu   hЏ @  �@���<EЏ^   hԨ<Ц�@4��	
Ԩ<Φ�@%Ԩ<��`� �@�P�������������������1���Ԩ��1��hЏb   �Ԩ<Џ�����@��ok ���1Ԩ<Ԩ@��Ԩ���X���A  1bЪ@��խ�*ѭ�p   ���P���c PV������@��fݏO� ���_  1� �
1� ѫ(ѫ)���P���P�@��j ��Э�P�@��j ��`���P��c �����P��c ����0 ݭ�ݭ�ݏj� ��,�  ���P� �c ѭ��Эح�Э�@ ֭��խ����P��c ݏz� ��9_  1� ѫ(?ѫ)9���P� �c ���P��c ݏ�� ��_  �fݏת ���^  U����ݏ�� ��\_  >��P�Pˏ�����Q�QP~Э�P�@��i ݭ����  �P�fݏ� ��^  �X��  �PX1��kЏa   P�Pk�PhЫ<Xˏ�����P�P ݏ3� ��\^  ��P�Pˏ�����Q�QP�Ы�Ы�1e�kP1� ݏG� ��%^  1oЏa   P�Pk�PhЫ<X��P�PP�PP� Pˏ�����Q�QP�Ы�Ы�15�� ݫ@���l����P��Џa   P�Pk�Phݭ�ݫ<�;��L����PX1� � Ы@Pݠ@���4����P��� Ы@Pݠ<�������P��Џa   P�P�@�Pk�Phݭ�ݭ���������Pݫ<��������PX1� ݏb� ��E]  1� �P�h   1�R�P;1F��P1 �
�P1���P1\���P�d   1���P�_   1����P�f   1����P�u   1���P�t   1��1s��P�v   1��1d�1a�1�ѫ�ݏ|� ��\  � �Z���#����PZ� �[�������P[Ъ��Ъ��Ъ��ݭ�ݭ�ݭ��Z�[ݏb   ��  �P[�Y$Џa   h�[X1k�h�[��n4  �P�<Ԩ@1Uѫ�ݏ�� ��\  1>ԭ�߭�ݨ@��u  �PZ�Z�@ѭ��J Э��J ˏ�����P�P ݏ�� ���[  ��P�Pˏ�����Q�QP�ˏ�����P�P�@   ݏū ��[  ��P�Pˏ�����Q�QP�Ы�Ы��k=ѻ<7Ы<Pՠ@.Ы<PѠ@� @   Ы<P��@Q��c ��ѭ�ѭ��hѨѨ	2�h��P�PP�PP� Pˏ�����Q�QP�� �X�������PX1#ݨ������P��ѭ�Э�P�P��P�1� �Yݏګ ��C[  1� �P�p   <�A�3�f���������������+��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������1�ӏ�   ���X��$  �PX�X��$  �P���1  �PX��z2 	�X��  Э�D�XP     ^Ь[ЬZЫY�k8&�Zݫ<�������P�<�Zݫ@�������P�@�[P1� �Y�� �Y�Y�[��Y  �P[ݫݫ�Y� �[ݏc   ���  �P[�Y�Y	� ݫ<�������P�<Џs   k� jP� P�PjP
� jP�PxPjݫݫ�Y������P���j�@���j�[���0      �    ^ЬZЬYЬ[��) �Y�Z�ZP��c ݏ� ��#�  �YX�ZP��c ݏ�� ��[X  1� �H�ac W1� �W�p  ݏ� ��X  �P1� �WZ�P1� �WP��c Ps�[t���! b�WP��c �WP2�c P�P�@��b �Z��1����P7�WP��c $�P9�ZP��c �WP��c ݏ.� ���X  �P�P�����X1?��P   �   ^Ь[ѫѫ�P�P�PVѫѫ�P�P�P���kXˏ����H�H PЫ<ZЫ@Y!Ы<Z�ZY�[P1��P�� ��   ���V�P�P�jP�[P1��V�P�P�iP�[P1��VPЩ<��Ѫ@� @  ѩ@� @  �[P1�ѩ@� @  �X�[P1�Ѫ@� @  �X�X�[P1l�H�SG �[P1Z�XP1t�V`��1����<Ѫ@� @  
Щ@�@Щ�1��Vb��­��<1��Vd��ĭ��<1��V q��/ ݏQ� ��V  f��1խ�ݏ_� ���U  խ�ݭ�ݪ<����  �P�<ƭ��<1�խ�ݏm� ���U  +խ�ݭ�ݪ<����  �P�<ǭ��<Pĭ�P�P�<P�P�<1?ҭ�P�P�<14ȭ��<1,̭��<1$Э�WxW�<�<1Э�W�W ݏ{� ��[U  1�խ��W P�WP�<�<�W P�WP�<�<1��Vr��Ϊ<�<1�Ҫ<�<1�ѪѪ�js��P�P�P�<ժ<�P�P�P�<1�Ѫ<���P�P�P�<1zѪ<���P�P�P�<1eѪ<���P�P�P�<1PѪ<���P�P�P�<1;í��<P�P�P�P�<1%í��<P�P�P�P�<1í��<P�P�P�P�<1� í��<P�P�P�P�<1� Ѫ<���P�P�P�<1� Ѫ<���P�P�P�<1� �[P1� �P�S   ����������������l�����w����������������������������������������������������������������������������������������*���������������������������������������1��[�F���p�����1G��ZYЏa   iݫݫݫ�Z��`  �PZЏa   k�ZP �   ^Ь[Ы<ZЫ@YЪXЩW�X
�W
.�X
�W

Ѫ�1��kP�@�A ݏ�� ��
T  1�ˏ����XP�P ˏ����XP�P�`   �YZЫ<Yˏ�����P�P Iˏ�����P�P�`   7�j ժ<Ѫ@� @  Щ�Щ�Щ��[ݏ�� ��  1ЪVЩ���XWѪ��[ݏ�� ���   1� ˏ����XP�P�`   ˏ����XP�P 1� ˏ����WP�P�`   ˏ����WP�P 1� ˏ����XP�P�`   5ˏ����WP�P�`   $Э�P�F��\ @��\ �[ݏϬ ��j   eˏ����XP�P�`   �Vˏ����WP�P�`   ֭�+�XP�Pˏ����XQ�QPX�WP�Pˏ����WQ�QPW1��[ݏڬ ��       d   ^мP�@��? ݬݏ� ߭���E�  ��� ߭���;R  
߭����P    �   ^Ь[Ы@P��@Q���c Q��Э�P��t �Џa   �@Џa   kݫ<��D  �P[ˏ�����P�P �)�Э�P��Q�QQ�QQ� QЭ�Pˏ�����R�RQZЭ�P2�YЭ�P2�X�X�Y�Z�[��  �P[Э�PР��Э�P��Wӏ@   W[Э�PРP'�V�X?�V�X7� V�X/ݏ � ��P   �P����������������������������V��P�VP��խ�/�X�Y�Z�X�Y�Zݭ���j&  �P�[���q  �P���'  �P[� �[���<����P[ӏ@   WGЭ�P2�~� Э�Pݠ� �[ݏg   ��*  �P[Э�P�V�Q�VQ�Q�QxQQˏ����WP�PQ�@�[��'  �P[�[P         ^Ь[�kP8Ы<[�ˏ�����P�P�`   ˏ�����P�P�@   �Pi�Pe�P`�P�u   �/�P�g   ��P��P���P�^   ���P�t   ���P�w   ��P�v   ���P�x   1r���      ^�� �� � ���(  �P[Ь�<Џ @  �@�[��&        ^Ь[ݫݫݫ�[��   �P���$         ^Ь[ˏ�����P�P ݏ� ��N  � P%ݫݫ��P�Pˏ�����Q�QP~�����       ^Ь[ЬZ�� ��[���  �P[�Z��T����P�[�<��7����P���%  �P[�� ��[��         ^Ь[ЬZ�Z�   Ы<Yݫ@�� ����PXЫ@Yݫ<�������PX�� ��Y��[  �PY�X�Y�������P��Z%  �PX�Z�   �X�<�X�@�[P        ^Ь[ˏ�����Z�Z
�ZkЫP�@��W �Z)ЫP�@��W  �ZЫP�@��W �Z�Z�Z��_����PZ�Z���P�ZP��k�Z�P�P��P�     ^Ь[ˏ�����P�P�`   )��P�Pˏ�����Q�QP�֫� �[�������sˏ�����P�P�@   � �[������Rݫ������PZ�Z��[P:�k�h   �[���   �P�ZP�P��P��Z� �Z�[���  �P[�[P       ^ЬPD�P1� �P1� � P1� � P1� �!P~�"Pyݏ*� ��zK  �Phݏ[� ��iK  �PW�P������������������ ����������ˏ�����P�P ˏ�����P�P�`   � Pݬݏ�� ��K        ^Ь[�k�h   ݏ�� ��iK  ѫѫ	ѫݏ�� ���J  �P)ݫ������PZЫ<Pݠ�������ZP�P�P      ^Ь[�kP}Ы<PРZ�Z�Zˏ����ZP�P ˏ����ZP�P�`   �k3Ы@PРZ�Z�Zˏ����ZP�P ˏ����ZP�P�`   �k�[P1� ݫ<�[��4���1� �P�Q   ��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����{�{�{�{����������kݏ˭ ���I  �[P �   ^Ь[�kWЫ<PРZ�ZXЫ@PРYЫ<PР��Ы@PРVЫ<PР��Ы@PР���WP1� 1� ݫ<�������P��ݫ@�����ѭ�Pݏ� ���H  �P�P��P�ԫ�[���   1� �ZYݏ�� ��H  1� ˏ����ZP�P �YX�V��Э���gˏ����YP�P Xݭ��Y�������P��ݭ��X������ѭ�P�YXЭ���,�P1H��P��P$18��P:10��P�r   1$�1~�ݭ�ݭ��Xݫ<��3  �P�<ݭ�ݭ��Xݫ@��  �P�@�G�8 �X�Э��Э���[��     �   ^Ь[�kZЫ<WЧYЫ@VЦX�fAѦ@� @  7�Y�Y
�Y�Y#�Yݦ<���  Ѧ<P�YX�X�Ч�Ч��gAѧ@� @  7�X�X
�X�X#�Xݧ<��  ѧ<P�XY�Y�Ц�Ц��Y�X�Z�r   ݏ� ��G  ԭ��Y�Y����
Y�X�X����
X�Y
�Y�X
�X�Y�X���T�Y�X���D�Y�X���4�Y�X���$�Y�X����Y�X�������Z:�Z�r   �Z$F�Y���Z$ѭ����ѭ�ѭ����Э�Y�Y��ѧѧ���ԭ�ЦXխ�"ѭ�ѭ�ӏ    J�6 �
����@ӏ    J�6 -����
YP�YP�P���X�X�Y	�Y�X��Э���ѭ�Yݭ�� ݭ��W��   �P�<ѭ�Xݭ�� ݭ��V��   �P�@�J�16 Э��ԫЭ���J�6 Bѻ<�h   8Ы<PР<WЧ��խ�ѭ�
ѭ��
��Э�P�P��P�Ч�Ч���� &ݭ��X�J�3 �Y�[ݏ5� ���  �[��  �[P   �    ^Ь[ЬZЬYЬXЫW�W
�k�[�����ЫWˏ����WP�P�`   ˏ����WP�P�@   �[��	����P[ЫW�ZW�kѫ@� @  �Z��Y��X��[P1� ӏ`   Z2ˏ����WP�P �k�b   ��X�Y�Z� �[ݏh   ���   1� �kCѫ@� @  9�Z�Z�k�W�Wn�<�n�<�1~��Zݫ<��  �P�<1k��W[�ZV�kPˏ����@�x4 Q�QA�kP�@�g4 4�k�F   +�X�Y�Zݫ<������P�<�X�Y�Zݫ@������P�@1��X�Y�Z� �[ݏh   ��            ^� �E  �P[ЬkЬ�<Ь�@Ь�ԫDЬ�Ь��[P         ^Ь[�kݏT� ���B  �ZЫ<Z�Z�<ݏn� ���B  �[��hE  �ZP   �    ^Ь[�Z�kWˏ����G�n3 P-Ы@Pݠ��  �PX�XZЫ<Pݠ��q  �PY�YP�PZ�P��
 
 
 ���WP1,Џ   P1E�Y�P1:1�Y�P1,1Џ  P1�P1�P1�Z� P1	1��Z� P1�1�� Y� X
Џ  P1��Z
Џ�   P1��Z
Џ�  P1��Z
Џ�  P1�1�Џ  P1�Џ   P1�� Z
Џ  P1��Z� P1��Z
Џ  P1w�Y�X�
P1g�Y�X�P1W�Z
Џ  P1H1,�Z
ЏE  P16�W�r   
�Y�$P1#�Z
Џd   P1� Y� X
ЏG  P1 �Z1��Y
ЏB  P1��Z
Џf   P1��Zݏ�� ���@  �P1�1��Z
Џ`   P1�1��Z
Џ`   P1�1��Z
Џ`   P1��Y�X
ЏD  P1y1]�Z
Џ�  P1g�X1F�Z� P1T�Y�X
Џ  P1@�Y�X
Џ  P1,1�P1#�P��   �����������������[����m����m��m�g�{���������g��[��m��m��m�q����������#�#�#�#�#�#���������������������������G��- ݏ�� ��?  �P        ^Ь[�[P"�PD�P?�P:�P5�P0�P+�P&�P���������������������������������      ^Ь[ЬZ�ZPTӏ�   [
ɏ ���[Paˏ ���[PWӏ �  [
ɏ  ��[PDˏ  ��[P:ӏ   �[� [P+� [P%�[P �P���������������������������      ^Ь[ݫݫݫ��K����PZ�[��@  �Zݏ̮ ��!?  �Z��T����P[���[P          ^ݏݮ ��n�  ݏ� ݬ��   ݏ� ��Q�       ^Ь[�kPˏ����@�L. Z�Z��d ݏ�� ݫ@��������N ��H Y�Yݏ�� ����  �Y��Yݏ�� ����  �kP�@��+ Ï [PǏH   P~ݬݏ�� ���  �Z ݫ<ݏ
� ���  ݫ@ݏ� ���  ݏ� ���  ݫ��5   ݫݫݏ%� ��j�  �Z�� ݏ7� ݫ<��������      ^Ь[ˏ����[P�P ݏ�� ��!�  Vˏ����[P�P�@   ݏ�� ���  6ˏ����[P�P�`   ݏ�� ���  �K� ݏ�� ��˿  �[P�Pˏ����[Q�QP[1w�      ^Ь[�[Y�Y�I�h; �Y��Y�_ �YP+��_ Z�Y�[Y�I�<; �  �Y�_ �ZP      ^Ь[�kZ������ЫY�Y� ~� ~��)�  � �b   �PZ�Z��N�  �Y	Џ@   ~� ~p�~��~  ԫ<�Z�@�k�kPˏ����@��+ Z�Z
ݫ@��u����Z
ݫ<��f���       ^��1 ��+ P         ^Ь[ЫD�^ �� 	�[��������� ݏ�� ���;  ��r� �[���  �P[�[��i  �P[�[������� ������[��   �[��
=        ^Ь[�� � �68  �[��   �[��H/     �    ^Ь[�kXˏ����H��* Zԫݫ�  �P��XP1� ѫ@� @  ԫ4|ի@$��@P��c ��R�  �PW�W���<  �P�4S��] Pѫ@P$Ϋ@~ݏȯ ߭���׿  ߭���<  �P�4"Ϋ@~ݏ̯ ߭��ﳿ  ߭���m<  �P�41� Ы<Yݩݩ�����P�4ݩ���׸���P�81� ݫݫ@�  ԫ4~�P�d   �F�P�_   1��P1�
�P1���P�^   ���P�c   ���P�b   1u���P�t   1���P�f   1Y���P�u   1���1}��Z
ݫ<��u����Z
ݫ@��f���      ^Ь[ЬZ�Z�kPR�Z�<�[PYݫݫݫ�Z�������P�[������8Ы@Y�i��Z�<�[P$Ы@Y�i��Z�<�[P�P�����������     ^Ь[ЬZ�kP&�ZP�P�<�P7�Zݫ<��U����P�<�P"�P�P��P��P�t   ��P�u   ��      ^ݬݬ�������P[ݬ���!����PZ�[ �P#�[�P�[ �P�[�P�P     ^��� (Ï �PǏH   P~ݏ� ���  ݬ��_���ЬPР��ˏ������P�P ˏ������P�P�`   �P1ԭ�мP1_��u ݏ� �  ݬ�����ЬPР@��Э�Pݠ������P[ЬPݠ�� ����[Piݭ�� ݭ�ݭ��������P��ݭ���#���ݭ���E  �P[ЬP�[�@��� (Ï �PǏH   P~ݏ
� ���  ݬ��v������Ѽ;Э�P19ЬPР<��Э�Pݠ��n����P[ЬPݠ��]����[Piݭ�� ݭ�ݭ���"����P��ݭ������ݭ���  �P[ЬP�[�<��Q (Ï �PǏH   P~ݏ(� ��a�  ݬ���������Э�P1� �P�G   ��� ��� [�� � � ��� � ��� ��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � � [��P    �    ^Ь[��i &Ï [PǏH   P~ݏF� ��z�  �[�������k�h   ݏ\� ��/5  Ы<XЫZШY�hW�W �Z�Z1� �hj��<Џ @  �@1� �W�h   %�X��]����PШ<�<Џa   h�[������1Z��ZY�Z�Z1� �Z�Z�Z
�Y�Y�[P1� �Z�Z�
Z�Y�Y�
Yˏ����YP�P �Y�ZY:ˏ����YP�P ˏ����YP�P�`   �[P1� �WEݫݨ<�������P�<Ы�Ы�Ы�Џa   k�X��"����P�X��A  �PX�XP^�[��h����P�[PL�W�h   1���W�W�W�t   	�W�u    �W�^   �G��# 	�W�g   �[P1n�       ^Ь[Ы<Zˏ�����P�P �[��0  K�� ��Z������PZ�j�h   �Z�������PZЫ�Ы�Ы�Џa   k�Z[�[���
          ^Ь[�k8!ݫ<�������P�<ݫ@�������P�@�[P+ˏ�����P�P � �[��������P[��[��    �   ^Ь[�� ݏe� ��ε  �[��A���ˏ�������ѭ�
ѭ�	�[�������kWˏ����G�" PЫ@YЫ<Z�[P1��P�� ��   ���[��-����PX�X[�X��h���1u�� ݏx� ��@�  �[������WP1~ѫ�#Щ���� ݏ�� ���  �[������[P1!ˏ�����P�P �[��"���	�[��3���1�Ъ���j�h   Hѭ�Bѭ�<�W=7�W?2Ъ<�<Џa   jЪ<Zݫݫݫ�Y������PY�Y������P�@�Y��9  �P1�թ<)�W!�W	�W�W�W�A   	�W�C   1tѩ<�W�W=1aݩ<��  �PV�WЏA   P�Pk�PW�V�<1(�Y���  �Pթ<11!�Y������P�@1 �jPyЏa   jЪ<Z#1� ݫݫ��O����P1� ���S �@�jЫ�Ы�Ы�Џa   k��d ݏ�� �  �Z�������ZP1�ݏ�� ��=0  W�P��P1z��P�F   1{��P�H   1o��P�_   1c��P�t   1W��P�u   1K��P�v   1B��1(ݪݪ������P��ѭ�R�[Z��P�Pˏ�����Q�QP�� �Z�������P[�W�d   	ЏF   jЏH   jЭ�P�P��P�Ԫ1�ѫѫ	+Џa   k��X ݏ�� ��y�  �Z�������ZP1��j к<Pӏ   @�m Џa   jЪ<Z1���j1X�j1���Y���  �P1BΩ<�<�P�Pk�PW�Wi�Z���  �P
�j�i�ZX�YP�P�<�PZ�XP�P�@�PY�W@�j;�i6ݪ@��  �P(Ъ<�<Џa   jЪ@Z��<�<Џa   j�[�����1��W$�j�Y��J  �PѺ@Ъ@P��<�<1� �W@�j;�i6ݪ@��  �P(Ъ<�<Џa   jЪ@Zª<�<Џa   j�[��F���1S�W2�j-�i(к<PЪ<P��<�<?�P��P�t   ��P�u   ��W1� �Y��  �P�ݩ<��]  �PVx�Vcݫݫݫ�Z��:����PZЏa   iЏa   k�Z������PZ��o &Ï [PǏH   P~ݏ�� �  �Z�������ZP1�Џ@   P�Pk�PW�V�<�W �Y��  �Pթ<Ω<�<�P�Pk�PW�Y���  �Pթ<�W�W1H�14�Y���  �P	ѩ<1/�1�j,�i'ÏP   kP2@� k�ZX�YP�P�<�PZ�XP�P�@�PY1�ݫݫ��K����P���P1� ˏ�����P�P /� �Y�������PYЭ�P�P��P�ԩ�Y������PY�Y�@� �Z���Q����PZЭ�P�P��P�Ԫ�Z��^����PZ�Z�<Э�P�P��P�ԫ�:k�[P1Oݫݫ������P���Pcˏ�����P�P /� �Z��������PZЭ�P�P��P�Ԫ�Z�������PZ�Z�<ѭ��P�P�P��P�ԫЏs   k�[P1� 1� �P�b   ����t���� ����
���������������� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � z������ ����������� � � � � ��� � � � � � ��������������������� � � � � � � � ��|���� ��� ���[P         ^Ь[�kPˏ����@�� Q�QPݫ@�������P�@ݫ<�������P�<�P��
 
 
 ���[�����        ^Ь[�[	�[P�P[	Џ����P�Z�[	�[[�Z��ZP         ^Ь[�kѫ@� @  ˏ�����P�P �P�P      ^� ������P[���<�P�P��P��[P       ^��a� ���L ��           ^�
ݏ� ���>�  ݏ� ��q)  ݏ�� ���  ����          ^ݏ&� ��B)  ݏ|�  ���ˮ        ^ݏ<�  �
�ﰮ  ݏ<�  ��  ݏ|�  ��  ����ݏ�� �  ݬݬ��d|���P��� ��  Э�P         ^�� �l� � ���$         ^Ь[� ��)  �PZ(�H kj�jPˏ����@�� Q�QPݫ@�������P�@ݫ<������P�<�P��
 
 
 ���ZP      ^Ѽ.ЬPР<[�k!Ы<Z�j�jѻ@Ы@YЫ<�@�Y�<ЬP       ^Ѭ2Ѭ,ˏ�����P�P ѬѬѬѬѬ7��q� .��h� �W ��]� ��W� � ��J� � �PHѬ>��4� 5��*� ��$� �OW ��� ��� �R ��� �E �P�P          ^ЬP
� P.�P)�P��P��P
��P��P��P��P�M   ��       ^��-� 
ݬ��c�    �    ^Ь[���P�PP�PP�[Pë`X�X1� �	�P�XP�Ѭ�� �����PVիЫP� ������PW�W�V�Xݫݬ��  �ZЫY�Z�L�ZZP�PP�PP�[P�Y`-�ZZP�PP�PP�[Pݠ��  �ZP�Z�PP�PP�PP�[P�`Y	�W��  �Y�� �����ի�W�  	�W��_�  1� ѬQիЫP� �L����PW�W�6 �ݬ�[��l   ݬ���(  ի�W��.�  	�W���  B�Z�Z�*�ZZP�PP�PP�[Pݠ�ZZP�PP�PP�[P�`���  �Z�ի
ݫ��ߊ         ^Ь[ݬ��i   �PZ���P�PP�PP��8� P�ZZQ�QQ�QQ�[Q}a`�Zx�~�Z~�[������Z�$���P�P~�Z�~�ZZP�PP�PP�P[~�����      ^�Z�ZP�P��ZZ��ZP�PY�YP�P[�Y�P�P[�Y�P�[P�[P       ^Ѭ�1� ���P�PP�PP��<� ���P�PP�PP��8� ���   ���P�P��� �ｉ  m���P�P�P�� �����P��ݭ����   ��p ��   ݬx�~��f������P�P�P�ݭ���F�  ݬ���P�P~��:���       ^ݬݬݏ;� �� �  ݬݏP� ����  Ь          ^� ݬݏV� ��ł        ^ݬݬݏf� �拓           ^ݬݏ� �          ^լx�~ݏ�� ��f�  x�P�P��R        ^ݬ� ��           ^ݬЬPݠ<��          ^��є �P�P ݏ�� ��"  ì PxP�Pì Q�倫 Q�Q R�QRPP�P �� ���^R �  ��{� ��P�  ��j� ��d� �c�        ^Ѭ�@   p���p��~ݭ�ݭ�ݏ�� ��q�  v���V��~ݭ�ݏű ��V�  ����Q       ^��%�  ��+E ��%E �  ��� P�@�� ��E ݏڱ ��	�  �� ��խ� ��� �����ݭ����D ݏ� ��ڀ  ��w ��q �(� � ������P���         ^��D ݏ�� �  ��D ݏ� �  � �����P�_�  ��c \� �����P[�[ݏ � ��V�  ݏ/� ��I�  ݏ=� ��<�  ݏE� ��/�  �[ݏP� �� �  ݏ^� ���  ��%c fݏf� ���  ��� ��� ݏ�� ���  ݏ�� ���  ��� ݏղ ���  ��я PxP~��Ə ݏ� ��y�  ��~C P���c P~��  �[�[�9�K�P���c Pޭ�Q(`a�	���K�*O ���K�M ��߭���  �[�     ^Ь[���k��Ȅ  �Pݏ�� ��!  �k�ﰄ  �Pݏ� ��	       ^��P� P��x��P�P~� �����P��B �Pݏ� ���~        ^��P���c P[����
2�~2�~ݫ������P����7��	ݭ�ݫݏ� ��|~  ݭ��k���  �Pݏ)� ��_~  0��ݭ��k���  �Pݏ9� ��<~  ݏH� ���       ^ЬPp���խ�ЬP��ЬP��      ^ݏf� ��         ^ݏu� ��~        ^Ь[�[ݏ�� ��^  � �  �PZ(�H kj� �  �PY(�H ki�:j�[�@�Y�<Џx   iԩ@�ZP         ^� �Ѕ  �Y�[�[�1� �K�Z�j-1� �Z�j1� ��R` �jPT�Z�j���?` �Zv��M �P�P�P�M ���  ���  ��` ��� F�j~ݏ³ ��  4�P�X   �������������������������������������������1a��Y�[1A�� �Y   �YP         ^Ь[�[� �x  �P[�kԫ4ԫ<��� �a  �PZЫ��[�<Џl   jЬ�4�ZP         ^ЬZЬYЬ[�[ݏѳ ���  �Yݏ׳ ��  � �  �PX�Z	Џn   PЏp   P�PhЫ��[�<�Y�4�Z�8�Z�kP�@� �k�kЏo   k�XP        ^Ь[ݫ<��  �P/ݫ@��K  Џa   kݏ����ݏ�����ݫ<��  �P[1� ݫ<��  �P�;kݏ����ݏ������[��  �P[b� �N����P��ݏ����ݭ��	ݫ<��e  �PYݏ����ݏ�����ݫ@��J  �PZЏa   k�Z�Y��  �P[ݭ��[��F����P[�[P      ^Ь[ݫ<���  �P/ݫ@��k  Џa   kݏ����ݏ�����ݫ<���  �P[1� ݫ<��   �P�;kݏ����ݏ������[��  �P[b� �n����P��Џa   kݭ�ݏ�����	ݫ<��~  �PYݏ����ݏ�����ݫ@��c  �PZ�Z�Y��  �P[ݭ��[��f����P[�[P       ^Ь[�kZ�ZP1� ի<ի4�P�P1� ݫ@������1� ݫ<������Pݫ@������P�P�P1� ݫ<������Pݫ@������P�P�P1� ݫ<��   1� Ы@Yݫ<��b����Pݩ<��T���vݫ<��p   �Pݩ@��:���\ݩ<��.����Pݩ@�� ����P�P�P7�P3�P1��P��P11��P1O��P;1��P�L   1a��        ^Ь[�kZ�ZP1� ի<
ի4�P�P1� ݫ@������1� ݫ<������Pݫ@������P�P�P1� ݫ<������Pݫ@������P�P�P1� ݫ<��K���1� Ы@Yݫ<��:����Pݩ<��T���vݫ<��H����Pݩ@��:���\ݩ<��.����Pݩ@�� ����P�P�P7�P3�P1��P��P11��P1O��P;1��P�L   1a��        ^Ь[�k;ݏ޳ ��)  ի<
ի@�[PЏa   kի<Ы@PЫ<P       ^Ь[ЬZ� �<  �PY�[�ZP�Z�[P�;iЪ��[�<�Z�@�YP       ^Ь[ЬZݏ����ݏ������[��8   �PY�Z�YP*�Y� ��  �PY�iԩ<ԩ4���Y�Z� ��t���  �   ^Ь[ЬZЬYЬX�kW�W�m   mЏa   P�Pk�P�@Ы@PР<��Ы<[�[������Pݭ��[��G���1��[��_����Pݏ�����[��(���1hݭ�ݏ�����	�[��q���1Qӏ   G� /ˏ����G�� P�P��:ݫ@��  �P�:�Z�Z$�Z�G�� �W�b   	�W�q   �Z�Z1� �G� 1� � �  �P�����Э�PԠ4Э�P��<Э�PЫ�� �z  �P��(�H ���Э�PԠ<� �`  �P�����Э�PЫ�Э�PЭ�<Э�PЭ�@� �6  �P���W�W��Э�PЫ�Э�P�[�<Э�PЭ��@Э�[�Z	1��W1Y� �����P��� �����P���;kЫ@��ݏ����ݏ�����ZЭ�Pݠ<������P��ݏ����ݏ�����ZЭ�Pݠ@�������P��Э�PЭ�@ݫ<������PCЏa   ��Э�Pݠ@��6  Э�@ݏ����ݏ�����ݫ<������P�<�[�����1x	ݫ<��w����PCЏa   ��ݭ����  Э�PР@�@ݏ����ݏ�����ݫ<��T����P�<�[��[���1'	խ�1� Э�Pՠ@@ݏ����ݏ�����Zݫ<������P��խ�
ݫ<��|  Џa   P�P���PkЭ�P1�ݏ����ݭ��	ݫ<�������P�<ݭ�Э�Pݠ@�������P�@Џa   ���[P1�Э�Pՠ@8ݭ�ݏ�����	ݫ<������P�<ݭ�ݭ�������P�@Џa   ���[P1Yݭ�ݏ�����	ݫ<��a����P�<ݭ���3����P��Э�Pݠ@��!����P��Э�PЭ�@ݭ�ݭ�� ������P��ݭ�ݭ���4����P��Э�PЭ�<�;��ݭ��[�����1��Zz�WP�Zp�P<5��l ��l l l l l l l ��l ����l ��l l l l l l l l l l l l l l l l l l l l l l ��l ��l ��l l l l l l ����l �����Z"�W�[��F���1B�W�[��U���11ˏ����G�� PX�ZЏa   k�P1Wݏ����ݏ�����Zݫ@������P�@ݏ����ݏ�����W;�~�Z~ݫ<�������P�<�P�� ��   ���Z�W;_ˏ����G�_ P>�;k�[�������P[�[P1��k�l   �[P1{Џa   kЫ<P1mЏa   k�P1a�P�� ��   ���[P1I�WP1��Y ÏP   WP�@�e�  P�Pk�PW�XYЏ����Xѻ@1� Ы@Pՠ<�Ы@Pՠ4��WPN�W�Y   	ЏQ   PЏP   P�Pk�PWл<P�@� 1� 8�X�[�����1��Y�[��q���1��P�P   	��������������������Џa   P�P�@�Pkݏ����ݏ�����ݫ<������P[�[�Y�W�������P[�X�[P1R�[�X� ������1Bݏ����ݏ�����ݫ<��G����P�<ݏ����ݏ�����ݫ@��+����P�@�[�Y�W������P[�X�[�X� ��v����P[�[P1�ݏ����ݏ�����ݫ<�������P�<�X�Y�	ݫ@�������P�@�[������1�Џa   k�Y�X�	ݫ<�����1��X	� �l����XP�P���Y	� �X����YP�PV�;kݫ<��7����P3ݏ����ݏ�����ݫ<��W����P�<�X�Y�	ݫ@��C����P�@1� ݫ@�������Pfݏ����ݏ�����ݫ@������P�@ի@/ݭ�ݏ�����	ݫ<�������P�<�Y�Y�	ݫ@�������P�@�X�Y�	ݫ<�������P�<-ݭ�ݏ�����	ݫ<������P�<�X�Y�	ݫ@������P�@�[������P���Xݭ�ݭ�������P���Y�Vݭ�������P��Э�P1A�X	� �#����XP�P���Y	� �����YP�PV�;kݫ<������P3ݏ����ݏ�����ݫ<������P�<�X�Y�	ݫ@�������P�@1� ݫ@�������Peݏ����ݏ�����ݫ@�������P�@ի@.ݏ�����V�	ݫ<������P�<�X�X�	ݫ@������P�@�X�Y�	ݫ<������P�<,ݏ�����V�	ݫ<��l����P�<�X�Y�	ݫ@��X����P�@�[��_����P[�Xݭ��[��X����P[�Y�V�[��F����P[�[P1 �X	� ������XP�P���Y	� ������YP�PV� �����P���Pݏ�����	ݫ<�������P�<Ы@��ݭ��V�ZЭ�Pݠ<������P��ݭ�ݭ��������P��Э�PЭ�<�X�Y�ZЭ�Pݠ@������P��Э�PЭ�@�;k�;���Y�V�[������P[�Xݭ��[��q����P[�[P1+ˏ����G��� P:ݏ����ݏ�����ݫ@��!����P�@ݏ����ݏ�����ݫ<������P�<�P��
 
 
 ���Y�[�YݏQ   ��L����P[�X�[�X�Y�~ЏP   ~��+����P[�[P1� �P�D   ��b��L�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b���b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b���b�b�b�J�J�J�J�J�J�J�J�J�J�1��     ^Ь[���z ݏ� իDЫD~��|. ~��p  ��z �[ݏ����ݏ������[�������P[�[�[��[  �[���  � ��s         ^Ь[ЬZ� [P� P�P[P
� [P�PxP[���  �.  �[�� ��. ��  ��� ���� �[��� �[���         ^� ��� P� P�P��� P� ��� P�PxP��� � �� P� P�P�z� P� �p� P�PxP�e� � �� P� P�P�� P� �� P�PxP�v� � ��n  ��i� ��c� �&� �� � �O�         ^ݬݏt� ݏ�B	 ��Mj  Џ�B	 P         ^Ь[��PR2�P�P�@�8 Z�Z.�J�, %�J�" P���c P~������P�P(�Z��P ���P�P�P
�������������      ^��59 ��~�4ݏ\� ��h          ^ݼ��n  �P��L  ݼ���m  �P��*, �$ݼݏ� ��@h  ݬ��         ^ݬ��        ^��8 :� ���  ���+ 	���+ ~���+ ~ݏ�   ݏ\� ���g  ��+      ^��+ P���c P[ݬ��e����Pݏx� ��g  ݏ�B	 ��}  ��+8 !ݏ�B	 ��Y+ ݏ�   �kݏ� ��lg           ^���7 �署 ݏ�   ݏ\� ��>g         ^���7 ��}� ݏ�   ݏ\� ��g         ^       ^Ь[��P4ˏ�����P�P�@   ��u7 �[������P	�[��5   $"�P����������    �� ��  ��        ^       ^Ь[ի1.��7 6��@�/ݫ��Pʏ����PxPPɫP~ݏp   �kݏ�� ��<f  1���P1ЫY�YP�YP�P~ݫݏ�   �kݏ�� ��f  1ݫݫݏ@   �kݏ�� ���e  1�ЫY�YP�YP�P~ݫݏ�   �kݏ�� ��e  1���P6 � ݫ� �kݏ�� ��e  1�ˏ�����P�P�@   � ݫ�2�kݏ�� ��qe  A��	ݫ������P~�k���j  �P~ݫ����
�(~�&~�kݏ� ��.e  13���5 1(� ݫݏ\   �kݏ�� ��e  2�P�P�@�1 X�X%�H�% �H� P���c P~��G����X�2�P�@�� ~ݫݏ^   �kݏ�� ��d  1^��=5 *ЫY�YP�YP�P~ݫݏ`   �kݏ�� ��ud  {��	5 ݫݫݏ`   �kݏ�� ��Pd  11ݫ�k��~ݏ|� ݏ�� �  ݏ�� ��}�  1� �P��`����`�����s�3���s������������ˏ�����P7��4 -� � ݏ�   2�P�P�@� Q��c ݏ�� ��c  
�P��������B4 YЫZ2�Xӏ`   ZHˏ����ZP�P�`   !�XP�X�@�� � ݏ�   ݏ,� ��_c  �ZP�Pˏ����ZQ�QPZ�     ^Ь[Џ�C	 Y��Z�Z"�Z��Z�Џ�C	 P         ^ݏ� ݏdC	 ���  �P�P1� ݏ� ݏdC	 ��(�  � �������P����5 eլ#� ������P��j����P��Pݏ�� ��b  ݬ��v& 	��n& ~��a& ~����  ݏdC	 ��-����Pݏ� ��fb  ��<& ���  �d   H� ��N�  �P����  ݏ�   ݏ� ݏ�� ��)b  ݏ� ݏ C	 ��^�  Џ�   �O�  խ�
ݭ��� ����P        ^��=� b� �������PU��l2 M� �������P����% 	��% ~��% ~ݏD   ݏ\� ��a  ��l% խ�
ݭ������    ^��D 1� ��yq ~ݏ�� ��Wa  ��eq ݏǴ ��Da  ��Rq �Mq P�PP�P~ݏݴ ��$a  ��2q ݏ� ��a  ԭ�Э�P��dC	 Э�P��dC	 ~ݏ�� ���`  ֭��ݏ�� ���`  Џ�� [�[�[��c fի_ˏ�����P�P�@   M��P'��@��71 �[��p����P	�[������ �P���� ��    �� ��  ���ݏ�� ��R`  � �g����P�������Pݏ� ��3`  ݏ�B	 ���# ݏ�   ݏ C	 �������Pݏ� ��`        ^���# ݏ� ݏ\� ݏ�� ��<}           ^���  ݏu   �����ݬ ݬݬݬݬݬݬݬݏ�� �	��|  ݏc� ݏ�� ���|  ��^�  ݏe� ��   ݏ�� ��{  ��>�         ^ݏc   ��>������  +���  "ݏu� ݏ�� ��~|  ݏ�� ��m{  \ݏ�� ݏ�� ��\|  ݬݬݬݬݬݏ�� ��@|  ݏ�� ݏ�� ��-|  ݏ�� ��{  ݏ�� ��{  ����y         ^��}�  Vݏw   �����ݏ�� ݏ�� ���{  ݬݬݬݏ�� ��{  ݏ�� ݏ�� ��{  ݏ�� ��z         ^Џ [�[��� Џa   k��H   [�Џ �4n         ^��!n [�[��� 
��H   [ZЏ Z�k�a   �Z��m �[P�Z[�[��m �ݏ¼ ��T���        ^��y�  ;�ZЏ [�[��� �k�a   �Z��H   [��Z�Zݏ� ������ ����Џx� ��  ��tm         ^Ь[�[@�kPˏ����@�
� Q�QPݫ@������ݫ<�������P��
 
 
 ��Џa   k     ^Ь[�[��N�  �PZ�Z��l P�P�   U����  ����  �h� ݏ � ��I������l ����  &ݏ   ���{  �PYݏ� ������Y���  �[��l ���  Y�Y�  �ZP�P�{l �YP       ^Џl� [�k�kPЫ@�� �kP�[@��� �[�       ^��!? \ݬݏ�� ���  ݬ��Y   ��g�  �
P��`�  Q��Y�  �Paݏ�� �
��w  ݬ��/	  ݬ��e���ݬ��	  ݬ��O���       ^����  P����  �P� �  լݏ�� ��-  1AмP�@�s ��խ�ݼݏ�� ��  1���P��@� ݏ�� ���~  ���P��<� P1����P��<� ݏ�� ���~  1�ݏ�� ��~  1�ЬPݠ��  ЬPݠ<��7���ЬPݠ@��)���ݏ�� ��|~  1�ЬPݠ��  ЬPݠ<������ݏ�� ��P~  1dЬPݠ<������ЬPݠ@ݏ�� ��+~  1?ЬPݠ@ЬPݠ<ݏ�� ��~  1!ЬPǏ@   �@~ЬPǏ@   �@Qď@   Q�Q�@Q�Qݏ�� ���}  ЬPݠ<��g���ݏ�� ��}  1�ЬPݠ���  ЬP2�:P� P~ݏ�� ��}  ЬPݠ<��"���ЬPݠ@�����ݏ�� ��g}  1{ЬPݠ��n  ЬPݠ<������ݏ�� ��;}  1OЬPݠ��B  ЬPp�~ݏ�� ��}  1)ЬPݠ4ЬPР8Q�A�[q P��@� ݏ�� ���|  ЬPݠ<��y���ݏ�� ���|  1�ЬPݠ���  ЬPݠ4ݏ�� ��|  ЬPݠ<��9���ݏ�� ��|  1�ЬPݠ4ݏ�� ��u|  ݏ � ��h|  1|ЬPݠ��o  ЬPՠ4<ЬPՠ<ЬPݠ<ЬPݠ4ݏ� ��*|  ЬPݠ4ݏ� ��|  ЬPݠ<ݏ� ���{  1ЬPݠ��  ЬPݠ<ݏ� ���{  1�ЬPݠ���  ЬPՠ<ЬPݠ<ЬPݠ4ݏ� ��{  [ЬPՠ4ЬPݠ4ݏ"� ��{  <ЬPՠ@ЬP��@Q��c ݏ'� ��^{  ЬPΠ@~ݏ,� ��G{  1[ЬPݠ��N  ЬPݠ<ЬPݠ4ݏ2� ��{  1/ЬPݠ4ݏ:� ��{  1ЬPݠ��  ЬPݠ4ݏ?� ���z  ЬPݠ<��q���1�ЬPݠ@ЬPݠ<ݏC� ��z  1�ЬPݠ@ݏM� ��z  1�ЬPݠ@ЬPݠ<ݏT� ��~z  1�ЬPݠ4ЬPݠ@ݏ]� ��`z  ЬPݠ<������ݏe� ��Ez  1YЬPݠ4ݏh� ��.z  ЬPݠ<������ЬPݠ@�����ݏm� ��z  1ЬP2�:~ЬPݠ4ݏp� ���y  ЬPݠ<��x���ЬPݠ@��j���ݏx� ��y  1�ЬPݠ4ݏ{� ��y  ЬPݠ<��8���ݏ� ��y  1�ЬPݠ��  ЬPݠ<ЬPݠ@ݏ�� ��_y  1s�P��   1�1� �P�^   �N�P1�� �P1���P1N�1C��P1��18��P%1���P$1��1#��P�F   1>�1��P�g   1��,�P�c   1]��P�b   1��1���P�d   1��1���P�n   1���P�l   1��1���P�t   1��1���P��  1��f�P��   1��,�P��   1���P��   1.�1u��P��   1��1f��P��  1���P��  1w�1I��P��  1��1:��P��  1R��P��  1��1��P��  1,�1�1�     ^ЬP1� ݬݏ�� �����Џ�� ��1Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� Џ�� ��1� �P��   �B�P��P1x��P1X�1E��P�1=��P ��P�1.��P�@   1=�1��P�   � �P�   1O�1��P�   1T�1���P�   1q�1��1��ݭ�ݏ�� ��v        ^ԭ����P��@� ���P��8� QЭ�A��j ֭��      ^��5 ݏ�� ��Vv        ^��b ����Ʌ ����tb ��nb ��Ь�8� ݏ�� ���w  �PV��� ��� ݏ�� ��\  ��� 1ݭ������� ��\  Э��+b Э��b ݏ�� �����1� ݬ���c  �P��Џ� �� Џ � ��m ���4 ѽ�(���PxP~ݏ� ��!\  �?� � ݭ���y   �P���� ��ݏ� �������f ��` �K� ��y4 -ѽ�('ݭ�ݏ4� ��IQ  ݭ������ݏ9� ��2Q  � �\  Э��Ka Э��{�    P   ^Ь��мP1R?ݼݏ;� ��s[  ЬP1�?ЬPѰ*ݬ��M  �ݏ�� ��v  ��#ЬPѰ#ݬ��K  �Pݏ�� ��[v  ȏ   �����dЬPѰ(ЬPРPݠ��/C  �PЬPЬQСQС�ЬPѰ(ЬPРPݠ���B  �PЬPЬQСQС�ݬ� ݏ   ЬPݠ�������P���� ��Э�P1�>���P�PP�PQ�Q�ݬ� ݏ   ЬPݠ�������P���� ��1���1ЬPݠ��nB  �P[ЬPݠ��]B  �[PЬPݠ��B  �P��1� ЬPݠ��5B  �P[ЬPݠ��$B  �[P3�� ���ݬ��SC  �ݏ�� ���t  ݬ��A  �P��5�� ���ݬ�� C  �ݏ�� ���t  ЬPݠ��A  �P�����PxPP��� P~���PxPP��� P~ݭ�ݏJ� ��KY  ������ЬP1v=���P�PP�PQ�Q�ӏ   ���
Э���Э����G���Э���Э��3���Э��ݬݬ���>  �P��ݬݬ���>  �P���P�ݬݬ��>  �P��ЬPѰ0:� �QZ  �P��ЬPРPΠQ�Q~ݏY� ���PxPP��� P~��O  9���PxPP��� P~���PxPP��� P~ݬ��0@  �Pݏ]� ��9X  ��PxPP��� P~���PxPP��� P~��t  �P<��PxPP��� P~���PxPP��� P~ݬ���?  �Pݏm� ���W  1� ӏ   �n���PxPP��� P~���PxPP��� P~ݬ��?  �Pݏ}� ��W  ��PxPP��� P~���PxPP��� P~���s  �PЭ���1�I��PxPP��� P~���PxPP��� P~���PxPP��� P~ݬ��?  �Pݏ�� ��W  ��1;��ЬP19;ݬЬPݠ��,A  �P���� ��Э�P1;ЬP� �(��ѭ���   ݭ�ݏ�� ��]���ݬ� ݏ
   ЬPݠ������P�����PxPP��� P��ѭ�?�� ��Э�P1�:ݬݬ��[B  �P��ݭ�ݭ�ݏ�� ��PV  ��Eݏ�� ���PxPP��� P~��Mr  ����PxPP��� P~��XW  ���PxPP�(�� ��Qӏ   �@���P�PP�PQ�Q�~� � ЬPѰЬPРPР~ЬPР~��$����P�Э�P1�9��PxPP��� P~���PxPP��� P~��r  �PЭ�P1�9��;ݬ��=  �P,���PxPP��� P~ݬ��R=  �Pݏ�� ��?U  10� ��,��PxPP��� P~ݬ�� =  �Pݏ�� ��U  1� ݬ���<  �P[ЬPݠ��<  �[PTѼNѼ%H��PxPP��� P~���PxPP��� P~ݬ��<  �Pݬ��<  �Pݏ�� ��T  1� ��:ݬ���<  �P+���PxPP��� P~ݬ��k<  �Pݏ�� ��XT  J��PxPP��� P~���PxPP��� P~ݬ��0<  �Pݏ� ��T  ݬݭ���Y  �P���ЬP1=8ЬPѰiЬPѰ_ЬPݠ���;  �P[ЬPݠ��;  �[P;ЬPРPݠ��w;  �P%ЬPЬQСQС�ЬPЬQСQС�1� ЬPѰzЬPѰ0pЬPРPՠcЬPРPݠ��;  �PЬPРPѠ��   )ЬPРPݠ��n;  �P#ЬPРPѠ� �  ЬPЬQСQС�ݬ� ݏ   ЬPݠ��Y����P���� ��Э�P17���P�PP�PQ�Q�ݬ� ݏ   ЬPݠ������P���� ��U�?� ݏ   ЬPݠ�������P���� ��ѭ�?�� ��ޭ�P�`P1�6�ݬ���;  �ݏ�� ��m  ���PxPP��� P~���PxPP��� P~ݬ��:  �Pݏ� ��R  �������ЬP1F6ЬPѰ!OЬPݠ��X  �P=��ݬݬ���7  �P�ݬݬˏ�����P�P~ЬPݠ������P��ݬ� � ЬPݠ������P���� ��Э�P1�5ݬݬˏ�����P�P~ЬPݠ�������P���� ��Э�P1�5��,��<��Pˏo���P����������PxPP��� P�� 1�Э�P1X5ݬ� ݏ   ЬPݠ��k����P���� ��Э�P1,5��*���Э�����P�PP�PQ�Q�~ݬ��6  �P���PxPP��� P~���PxPP��� P~ݬ��8  �Pݏ&� ��P  ��ЬP1�4ЬPѰ1� ЬPРPѰ#1ݬݬ��@6  �P�ݬݬݏ   ЬPݠ������P��;ݬݬ��6  �P�����P�PP�PQ�Q�~ݭ�ݏ   ЬPݠ��]����P���� ��ЬPݠ��=  �ݏ�� ��k  ݬ� ݏ   ЬPݠ������P��ݬ��7  �P[ݬ��7  �[P��Э�P1�3�� ��Э�P1�3��-���ݬݭ�ݬ���O  �P�ݬݬ��85  �P�ЬPݠ��7  �Pkݬ��d7  �P[ЬPݠ��S7  �[PKݬ��7  �P�f   ݬ���6  �P�d   
Џ6� ��ݬ��X>  �ݏ�� ��j  Џ;� ��ݬ��u6  �P[ЬPݠ��d6  �[P1� ݬ���6  �P[ЬPݠ��6  �[P]ݬ��26  �Pm��PxPP��� P~���PxPP��� P~ݬ��F6  �Pݏ?� ��3N  ݬݭ����S  �P�1� ݬ��Q6  �P[ЬPݠ��@6  �[PJ��PxPP��� P~���PxPP��� P~ݬ���5  �Pݬ��5  �Pݭ�ݏN� ��M  J��PxPP��� P~���PxPP��� P~ݬ��5  �Pݏ^� ��|M  ݬݭ���S  �P���ЬP1�1Џ������Џm� ��ЬPѠ	ݏq� ������ЬPѰ*ݬ��e?  �ݏ�� ��Ph  ����P�PP�PQ�Q�~Ь~� ݏ    ЬPݠ��N����P���� ��Э�P11� � � ЬPݠ��'����P����1������P�PP�PQ�Q�~ݬ��2  �P���PxPP��� P~���PxPP��� P~ݬ��N4  �Pݏ�� ��WL  ��@ ��Fѭ�
Џ�� ��Џ�� �욭�PxPP��� P~ݬ��4  �Pݭ�ݏ�� ��L  <���PxPP��� P~���PxPP��� P~ݬ���3  �Pݭ�ݏ�� ���K  ��1� ��� �l��PxPP��� P~ݏ�� ��� ��9B  Ï� ��� PǏ   PQ�Q���   ��� �� �������� �H�  � �Z  ЬP1�/�� �i��PxPP��� P~ݏ�� ��� ���A  Ï� �� PǏ   PQ�Q���   �n� �������`� ���  � �Y  ЬP1/ݏ�� ��z����� �ЬP1/��@ ��Fѭ�
Џ�� ��Џ�� �욭�PxPP��� P~ݬ��s2  �Pݭ�ݏ�� ��yJ  <���PxPP��� P~���PxPP��� P~ݬ��52  �Pݭ�ݏ�� ��;J  ��Э���1��� ��Э�P1].ЬPѰ*ݬ��M<  �ݏ�� ��8e  ݬ��<8  �P1�(ȏ   �ЬPݠ��/2  �PЬPݠ��2  �PЏ�� ��1�Џ�� ��ЬPѰ#ݬ��F>  �P�ݏ�� ���d  ЬPݠ��1  �P/���ЬPР�����ݬ� �K  �P�߭�������P�� ݬ� ��J  �P�ЬPݠ������P���� ��Э�P1R-���P�PP�PQ�Q�ЬPݠ��61  �P/���ЬPР�����ݬ� �J  �P�߭���4����P�� ݬ� �hJ  �P�ЬPݠ������P���� ��U��ѭ�?/ݭ�� �5J  �P�ЬPݠ�������P���� ��Э�P1�,�ݬ���1  �ݏ�� ��c  ���1��ЬPѰ*ݬ��n:  �ݏ�� ��Yc  ȏ   �Џ�� ��ӏ   �(��#ЬPѰ#ݬ��t8  �Pݏ�� ��c  ݬ� ݏ   ЬPݠ��,����P���� ��Э�P1�+���P�PP�PQ�Q�ݬ� ݏ   ЬPݠ�������P���� ��x��ѭ�?,ݭ�� ݏ   ЬPݠ�������P���� ��Э�P1�+ӏ   �ЬPѰ#�ЬPݠ��0  �ݬ��0  �ݏ�� ��@b  ݬ�� /  �P[ݬ���.  �[P1Tݬݬ���,  �P�����PxPP��� P~���PxPP��� P~���PxPP��� P~ݬ��.  �Pݭ�ݏ � ��F  ��ӏ   �Э��Э��ݬ��%.  �P~ЬPݠ��.  �Plݬ��.  �P[ЬPݠ��p.  �[PL��PxPP��� P~���PxPP��� P~ݬ��	.  �Pݏ� ���E  ݬݭ���K  �P�E��PxPP��� P~���PxPP��� P~ݬ��-  �Pݬ��-  �Pݏ!� ��E  ��ЬP1�)��1)���ӏ   �1� Э�����a3��@ ��+���PxPP��� P~ݬ��2-  �Pݏ2� ��;E  v���s3��@ ��+���PxPP��� P~ݬ���,  �Pݏ>� ��E  <���PxPP��� P~���PxPP��� P~ݬ��,  �Pݭ�ݏJ� ���D  ��1p��)���PxPP��� P~ݬ��,  �PݏY� ��D  ��ЬP1�(���Э��ݬݬ��V*  �P���Nӏ   �D���PxPP��� P~���PxPP��� P~ݬ��,  �Pݭ�ݏf� ��D  Э���1`�ݼ���D  �P=��PxPP��� P~���PxPP��� P~��f`  �PЭ��Э���Ь��1L���PxPP��� P~���PxPP��� P~��)`  �P1���PxPP��� P~���PxPP��� P~���PxPP��� P~ݬ��D+  �Pݭ�ݏu� ��JC  ��1� ��� �Lݏ�� ��PxPP��� P~��<_  ���PxPP��� P~��GD  ��PxPP�(�� ЬP1)'�� �5���PxPP��� P~��D  ��PxPP�*�� �� �ЬP1�&�� �ЬP1�&��ЬP1�&ݬ� ݏ    ЬPݠ�������P���� ��Э�P1�&��ݬݬ��J(  �P��� ��yЬPѰ#oЬPݠ��r*  �P\��Ь��ݬݬ��(  �P�����PxPP��� P~���PxPP��� P~ݬ���)  �Pݏ�� ���A  Э�����PxPP��� P~���PxPP��� P~ЬPǏ@   �Qď@   Q�Q�Q�QЬPǏ@   �~ЬPݠ���)  �P	Џ�� ~Џ�� ~ݏ�� ��^A  ��ЬP1�%ЬPѰ#ݬ� ݏ   ЬPРPݠ������P��ݬ� ݏ   ЬPݠ��u����P��ЬPݠ ��C  �P����XЬPѰЬPРPѠݭ�ݏ�� ���@  ,ݭ욭�PxPP��� P~ݬ��(  �Pݏ�� ��@  hЬPѰ2ݭ욭�PxPP��� P~ЬPݠ��V(  �Pݏ�� ��_@  ,ݭ욭�PxPP��� P~ݬ��((  �Pݏ�� ��1@  ЬPݠݏ�� ��@  ����� ��E ��E PxP~ݏ�� ���?  Э�P1'$ݬݬݬЬPݠ��<����P��ЬPݠݏ� ��?  ��N ��BE ��;E PxP~ݏ
� ��?  Э�P1�#ݬݬˏ�����~ЬPݠ�������P����/���)���PxPP��� P~ݬ��/'  �Pݏ� ��8?  ЬPݠݏ)� ��$?  Э�P1Y#ЬPՠHЬPՠ#ЬPݠЬPݠݏ4� ��]� ��5  ЬPݠݏ:� ��A� ��n5  ЬPݠݏ=� ��%� ��R5  ������ ���?  �$�� ԭ�ЬPՠ!ЬPՠ� ��ЬPѠЏ@   ��ԭ���1����Ѽ0��HÏ� �� PǏ   PQ�Q����   �� ������������� ���  � �L  Э�P1@"ӏ   ��a���^� ��/?  �*�P� Ï� �E� PǏ   PQ�Q����   �-� �� ������������ ��  � �TL  Э�P1�!ӏ�   ��qݏ@� ���� ��Y  ����� ��>  �(��� Ï� ��� PǏ   PQ�Q����   �� ������������� ��  � ��K  Э�P1Z!��� ����   �w� ݬݬ���"  �P�����PxPP��� P~ݭ�ݬ���$  �PݏB� ���<  ��1���1� ݬ���$  �P��� ݏQ� ��<  cݬ���$  �P%��PxPP��� P~���� ݏ]� ��h<  /��PxPP��� P~��� ݬ��J$  �Pݏk� ��7<  1$� ��,��PxPP��� P~ݬ��$  �Pݏ{� ��<  1� ��PxPP��� P~��X� ݬ���#  �Pݏ�� ���;  �� �:�+��PxPP��� P~��.J  �P�-��PxPP��� P~��J  �Pӏ   ��&�+���� ���I  �P\�-���� ���I  �PIÏ� ��� PǏ   PQ�Q����   �� ������������� ��  � ��I  Э�P1R��  ���ЬP1A���Џ�� ��1��� � �ЬPݠ��J����P�����PxPP��� P~ݏ�� ���:  ЬP1�ݬ���"  �P
ݬ��u(  ݬ���(  �P1>ЬPѰ*ݬ��,  �ݏ�� ��U  ȏ   ���#ЬPѰ#ݬ���*  �Pݏ�� ��wU  ݬ��o"  �P
ݬ���'  ݬ� ݏ   ЬPݠ��s����P���� ��Э�P14���P�PP�PQ�Q�ݬ� ݏ   ЬPݠ��9����P���� ��1D� ��yЬPѰ#oЬPݠ���!  �P\��Ь��ݬݬ��s  �P�����PxPP��� P~���PxPP��� P~ݬ��=!  �Pݏ�� ��F9  Э�����(���
ӏ   �Э��ݬݬ��  �P�ݬ��F!  �P1� ݬݬ���  �P�����PxPP��� P~���PxPP��� P~���PxPP��� P~ݏ�� ��8  ��PxPP��� P~���PxPP��� P~ݬ��   �Pݏ�� ��{8  ӏ   �-���PxPP��� P~���PxPP��� P~ݏ�� ��D8  ��ЬP1uЬPѰ01� ЬPРPР��ѭ�곏� �ⳏ @��ښ�PxPP��� P~���PxPP��� P~��nT  �P@׭���PxPP��� P~���PxPP��� P~���PxPP��� P~ݏ�� ��7  Э�P׭��P/��PxPP��� P~��PxPP��� P~ݏ�� ��f7  �1� ӏ   �?���PxPP��� P~���PxPP��� P~���PxPP��� P~ݏ� ��7  =��PxPP��� P~���PxPP��� P~���PxPP��� P~ݏ� ���6  ӏ   �X���PxPP��� P~��PxPP��� P~��6S  �P-��PxPP��� P~���PxPP��� P~ݏ&� ��y6  ��ЬP1�ЬPѰ*ݬ��(  �ݏ�� ��Q  ݬ��$  �P1�ȏ   �Џ4� ��ݬ��\  �P^ЬPѰ0%ЬPРPՠЬPРP���ݬ��p  ЬPѰ0%ЬPРPՠЬPРP���ݬ��A  1��ЬPѰ*ݬ���'  �ݏ�� ���P  ݬ���#  �P14��#ЬPѰ#ݬ���%  �Pݏ�� ��P  ȏ   �ЬPݠ��  �PЬPݠ��  �PЏ8� ��1y�ݬ� ݏ   ЬPݠ��v����P���� ��Э�P17���P�PP�PQ�Q�ݬ� ݏ   ЬPݠ��<����P���� ��1G횭�P�PP�PQ�Q�ݬݬ��  �P�����PxPP��� P~���PxPP��� P~���PxPP��� P~ݬ��T  �Pݏ=� ��]4  ���PxPP��� P~���PxPP��� P~ݬ��  �PݏP� ��$4  ���PxPP��� P~���PxPP��� P~���PxPP��� P~ݬ���  �Pݏ`� ���3  ��1$�ӏ   �Э��1ި��Э�P1�ЬPѰ*ݬ���%  �ݏ�� ���N  ݬ���!  �P10ȏ   �Џs� ��1`�ЬPՠ,ЬPՠ#ЬPݠЬPݠݏw� ��� ���)  ]ЬPՠЬPݠݏ}� ��� ��)  8ЬPՠЬPݠݏ�� ��e� ���N  ݏ�� ��P� ��})  ԭ�Џ   ��1i�ЬPѰ*ݬ���$  �ݏ�� ���M  ȏ   �Џ�� ��1��ЬPѰ*ݬ���$  �ݏ�� ��M  ݬ��   �P1ȏ   �Џ�� ��1C�ЬPРQ�A���  ݏ�� ��� ���(  ԭ�Џ�   ��ЬPѠ���1���ݬ���  �P�������1J�Э�P1.ݬݬ���  1ЬPѰ*ݬ��$  �ݏ�� ���L  ݬ���  �P
ݬ��z  ݬ���  �P1Cȏ   �ЬPݠ��  �P
ݬ��D  ݬ� ݏ   ЬPݠ������P���� ��Э�P1�ЬPѰ0C�� ��ЬPѰ#ЬPݠ��V  �P�� @��1� ЬPݠ��8  �P곏 ��#ӏ   �ݬ��  �ݏ�� ��L  ӏ   ���Э�����P�PP�PQ�Q���Ь��ݬݬ��  �P�����PxPP��� P~���PxPP��� P~ݏ�� ��_0  Э������P�PP�PQ�Q���(ӏ   ����Э��ݬݬ��  �P�����P�PP�PQ�Q�ݬ��?  �Pݬݬ���  �P��ӏ   �Э���Ь��ЬPѰ0GЬPРPР��8���PxPP��� P~���PxPP��� P~í� ~ݭ�ݏ�� ��/  1��ݬ� ݏ   ЬPݠ�������P���� ��1�皭�P�PP�PQ�Q�~ݬ��3  �P���PxPP��� P~���PxPP��� P~ݏ�� ��/  ���PxPP��� P~���PxPP��� P~���PxPP��� P~���PxPP��� P~ݏ�� ���.  1�ЬPаP1%ݬ� �ЬPݠ��
����P�����PxPP��� P~ݏ�� ���� ��%  ԭ�Э���1
�ݬ� �ЬPݠ�������P�����PxPP��� P~ݏ�� ��� ���$  ԭ�Э���1��ݬ� �ЬPݠ��|����P����� ��3���PxPP��� P~ݏ�� ��X� ��$  �����Џ   ��1oﳏ ��.���PxPP��� P~ݏ�� ��� ��J$  �����ԭ�19ﰏ ��Э�P1��P,�e�����ЬPР��ѽ�
1� ӏ   �xЭ�PѰ0nЭ�PѰ-dݬ��  Э�QСQ�P�Lݬ� �Э�Pݠ������P�����PxPP��� P~ݏ�� ��s� ��#  Џ H  �������1��ѽ�1�Э�PѰ�ӏ   ��Э�PРPѰ0�ݬ���  Э�QСQСQ�P��ݬ� ݏ   Э�PРPݠ�������P���� ��Э�P1����P�PP�PQ�Q���� ��zݬݬ��F  �P�����PxPP��� P~���PxPP��� P~ݭ���  �Pݏ�� ��,  ���P�P����P�PP�PQ�Q�Э������ ���� ��Э�P1%ݬ� ݏ
   Э�Pݠ��8����P���� ���ݭ���<  �ݏ�� ���F  ���PxPP��� P~���PxPP��� P~ݏ� ���� ��"  Џ   �����P���Q�QP��1��ѽ�1Э�PѰ0�ݬ� ݏ   Э�Pݠ������P���� ��Э�P1[��� ��dݬݬ���  �P�����PxPP��� P~���PxPP��� P~ݭ����  �Pݏ	� ���*  Э������ ���� ��Э�P1����P�PP�PQ�Q�ݬ� ݏ   Э�Pݠ�������P�����PxPP��� P~���PxPP��� P~ݏ� ���� ���   Џ   �������1��ѽ�1� Э�PѰ0�ݬ� ݏ   Э�Pݠ������P���� ��Э�P1B��� ��dݬݬ���  �P�����PxPP��� P~���PxPP��� P~ݭ���  �Pݏ� ��)  Э������ ���� ��Э�P1����P�PP�PQ�Q����PxPP��� P~Э�PРPΠ~ݏ.� ���� ���  Џ   �������1��ѽ�1� ӏ (  �xЭ�PѰ0nЭ�PѰ-dݬ��X  Э�QСQ�P�Lݬ� �Э�Pݠ��a����P�����PxPP��� P~ݏ5� ��E� ��r  Џ H  �������1\�ѽ�dЭ�PѰ-Zӏ   �PЭ�PѰ-Fݬ���  �P7Э�PРPݠЭ�PРPݠݏ;� ���� ��  Џ   ��ԭ�1��ݬ� ݏ   ЬPݠ������P���� ��Э�P1h���P�PP�PQ�Q��� ��.���PxPP��� P~ݏF� ��f� ��  ԭ������1�鳏� ��eݬݬ���  �P�����PxPP��� P~���PxPP��� P~ݭ���  �PݏJ� ��'  ���P�P����P�PP�PQ�Q�Э������ ���� ��Э�P1����PxPP��� P~ݏY� ��� ���  ԭ������1��ЬP��$Q�Q1Џl   ��ݬ� ݏ
�  ЬPݠ��n����P���� ��Э�P1/���P�PP�PQ�Q�ݬ� ݏ
�  ЬPݠ��4����P���� ��U�?� ݏ
�  ЬPݠ������P���� ��ѭ�?�� ��ޭ�P�`P1�
�ݬ���  �ݏ�� ��A  ���PxPP��� P~���PxPP��� P~ݭ�ݏ^� ��;&  ӏ �  �ݭ�ݭ����)  �P��Э�P1U
ЬP��$Q�QЏq   ��1��Ѭ?�� ��Э�P1)
ݬ� ݏ�  ЬPݠ��<����P���� ��Cݬݬ��  �P�����PxPP��� P~���PxPP��� P~ݏm� ��%  Э������P�PP�PQ�Q�ݬ� ݏ�  ЬPݠ�������P���� ���ݬ���  �ݏ�� ��q@  �� ��Cݬݬ��  �P�����PxPP��� P~���PxPP��� P~ݏ{� ���$  Э���ݭ���'  �P���� ��6ЬPѰ#ݏ�� ������ЬPݠ��3  �ݏ�� ���?  ݭ���6'  �P���� ��6ЬPѰ#ݏ�� ����ЬPݠ���  �ݏ�� ��?  ���PxPP��� P~���PxPP��� P~ЬP��$~ݏ�� ��$  ӏ    �(�?ݬ���  �P��ЬP��$~ݏ�� ���#  ���Э�P11����Ѵ  ЬPݠݏ�� ��2� ��_  ԭ�Џ   ��1K��林  ЬPݠݏ�� ��� ��1  ԭ�Џ   ��1�ݬ� ݏ    ЬPݠ�������P���� ��Э�P1����P�PP�PQ�Q���ݬݬ��'	  �P���� ��Lݬ��  �P�����PxPP��� P~���PxPP��� P~ݬ���
  �Pݏ�� ���"  Э��������PxPP��� P~ݏ�� ��"  9��PxPP��� P~���PxPP��� P~ݬ��
  �Pݏ� ��"  ��w��� �Gݏ� ��PxPP��� P~��v>  ���PxPP��� P~��#  ��PxPP�(�� (���PxPP��� P~��W#  ��PxPP�*�� ЬP19ԭ�1B�ݬ� ݏ   ЬPݠ��F����P���� ��Э�P1��*���Э�����P�PP�PQ�Q�~ݬ��  �P���PxPP��� P~���PxPP��� P~ݬ��Z	  �Pݏ� ��c!  ��ЬP1�ԭ�1��ЬPѰ2=��8ݬݬӏ    �	Џ    P�P�P~ЬPݠ��~����P��Э�P1GЬPѰ3
ЬPѰ1dݬݬӏ    �	Џ    P�P�P~ЬPݠ��2����P���� ��Э�P1�Э���� � ݏ    ЬPݠ������P�1��ЬPѰ*1rݬ� ݏ   ЬPРPݠ�������P�����P�PP�PQ�Q�ЬPѰAݬЬPݠ��,  �P�����P�PP�PQ�Q�~ݭ�ݏ   ЬPݠ��z����P��ݬ� ݏ   ЬPݠ��[����P���� ��/�ЬPРPݠ��W	  �ݬ��K	  �ݏ�� ���:  �$�����PxPP��� P~ЬPРPǏ@   �Qď@   Q�Q�Q�Qݭ�ЬPРPǏ@   �~ݭ����PxPP��� P~ݏ.� ��Q  ��1��PxPP��� P~���PxPP��� P~ݏF� ��  ���Э�P1P��1VЬPѰ#��Ь��ݬݬ���  �P��ݬݭ�ݏ   ЬPݠ��2����P���� ��Э�P1����P�PP�PQ�Q�ݬ� ݏ    ЬPݠ�������P���� ��\��ѭ�?8ݭ�� ݏ    ЬPݠ�������P���� ��Э�P1�ݬ��_  
ݬ��{  �ݏ�� ��b9  ���PxPP��� P~���PxPP��� P~ݬ��  �PݏT� ���  ��PxPP��� P~���PxPP��� P~��T:  �P��ЬP1�1�ЬPѰ*Mݬ���  �P>ݬ���
  ݬ���  �P�P�P�P[ЬPРP�[��ݏ�� ��8  ݬ� ݏ    ЬPݠ������P�����P�PP�PQ�Q�ЬPѰ!
ݬ���  ݬݭ��ЬPݠ��r����P���� 4��1� �� ��O��ѭ�?)ݭ�ݭ��ЬPݠ��:����P���� ��Э�P1� ݬ���	  �ݏ�� ���7  1ӏ    �'������ݬ��  �ݏ�� ��7  ��Э���1����)<��Pˏo���P����������PxPP��� P醴 1��Э�Pm�P2���,�#����H����(�s������s���w��^�����K������0�K���˰���Bܟ�k��0�6���7���٪�N����|���;��1A�        ^��%� P��� �,P��hL P����� �   ݏX� �בּ��Э�P      ^ѼЬ����
ЬPРPЬPРP�P��� �����P��Э�PЭ�QС�ݭ���d  �P�P�P�P����R���P���C PD�-��Э�P���C Qí�Q�Э�P��­��C ����  �C ��C ��  Э�P�,��ݭ���y  �P[Э�P�[�Э�P         ^�  ݬ��  �P�~�~��7  �Pݏo� ��͵ ��*6  Ï� ﻵ PǏ   PQ�Q����    �������� ��  � ��(  Э�P         ^ЬPѠ
������ԭ�ѭ�1� x��P�P�1� ѭ��P�P���QxQQ�Q��Q�Q�QP1� Э�P�@�[�  ݏv� ��� ��0  x���ѭ����PxPP�P�Ï� �ش PǏ   PQ�Q����   ��� ��� �������ﯴ �&�  � ��'  Э�P1� ֭�18�� ݬ������P��ѽ�-hЭ�PРQ�Aﻩ  ݏy� ��c� ��  Ï� �Q� PǏ   PQ�Q����   �9� ��� �������*�   � �d'  Э�Pf�  Э�Pݠݏ|� ���� ��*  Ï� �� PǏ   PQ�Q����   �ӳ ���������ĳ �;�  � ��&  Э�P          ^ЬPѠ	
ЬPѠ
�P�P        ^ЬPݠ��            ^ЬPРP��� P        ^ЬPРQ�A�ب  P       ^ЬPРQ�A��  P       ^ЬPРQ�A��  P      ^� �����P��мP1� ЬPݠ�������P��ЬPݠ�������P��(,���Э�PЭ��Э�PЭ��Э�P1� ЬPݠ������P��(,���Э�PЭ��Э�P1� (,���Э�P{ݏ�� �����l�P2v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v�v����������������������������������������������       ^� �����P��ݬݬ�������P��� �����P����ЬP(,���
ЬP(,������Э�PЭ����Э�PЬQС�Э�PЬQС����Э�PЭ��Э�PЭ��Э�PЭ�QС���ЬPЭ��	ЬPЭ��        ^мP1yݬЬPݠ�������P��ݬЬPݠ�������P��Э�P1p� �$  �P��ݬݭ��ЬPݠ��ƹ���P��<��Pʏ����P1=Ѭ?
Џ   P1-ݬ� ݏ
�  ЬPݠ����P��ЬP��$��ЬPѰGѭ�Aѭ�;ݭ�ݏ�� ���  ݭ�ݏ�� ���  ЬP��$~ݏ�� ���  �P1� ѭ����PxPP��� P~ݏ�� ��  [ѭ����PxPP��� P~ݏ�� ��|  6ݭ�ݏ�� ��j  ���PxPP��� P~ЬP��$~ݏ�� ��D  <��Pʏ����P(�P��$ $ $ $ $ $ $ $ $ $ $ $ $ $ ��$ ��       ^ЬPѠ
�P�P�P�����ѭ�����  ݏ� ��9� ��f
  ҬP�P��ݏ� ��  Ï� �� PǏ   PQ�Q����   ��� ��� ���������� �^�  � �!"  Э�P        ^� �����P��(,���Э�PЬ����Э�PЬ�Э�P       ^� �\����P��(,���Э�PЬ����Э�PЬ�Э�P       ^� �$����P��(,������Э�PЬ�Э�PЬ�Э�P       ^� ݬ��+����P��ݭ�ЬPݠ��.����P��ЬPР��ѽ�,ݭ�ݭ�Э�Pݠ������P��n����P��Э�PР���ݭ�ݭ�ݭ�������P��F����P��(,���        ^� �\����P��� �Q����P���P�P���P��Э�P�QЭ�R�Q��Q�Э�PЬQС�Э�PЬQС�ЬPѰ0	ЬPЭ��ЬPЭ��     ^ЬPѰ�P1ЬPРPѰ#ݬ���  �Pݏ�� ��,  � �����P��(,���мP1� ���1� ���1� ���1� ���1� ЬPݠ�������P�P1� ���rЬPݠ�������P�P1� ���UЬPݠ������P�Ps���9ݏ*� ��
���*�P{������������������������������������� ������P��ЬPРP(,�����ЬPЭ��ЬPЭ���P       ^� �����P��(,���Э�P��ЬPЭ��    ^�ݏC� ���".  ЬPРPРPР��ЬPР��� ݭ�������P��� �I����P�����Э�PЬQС�� �-����P[Э�P�[�Э�P��Э�PРPЭ�QС�Э�PРPЭ��Э�PРPЭ��� ������P[Э�P�[�Э�P(,��ЬPРPРPЭ��(,��        ^� �����P�����Э�PЬQС�� �����P�����Э�PԠЭ�PЬQСQС�Э�PЭ��� ݭ�������P��Э�PԠЭ�PЭ��� �<����P�����Э�PЬQС�� � ����P��(,���Э�PЭ�Э�PЭ��Э�PЭ�QС�Э�PРPЭ��(,����P        ^� ������P�����Э�PЬQС�� �����P�����Э�PԠЭ�PЬQСQСQС��ݭ��������P��Э�PЭ��� �l����P��(,���ֽ�Э�PРPРPЭ��� �G����P��(,���Э�PЭ�Э�PЬQСQС����(,���ЬPЭ��ЬPЭ��P      ^ЬPРPР��ѽ�#ݬ���   1� Э�PР��� ݭ�������P��� �����P��Э�PЭ�QС����Э�PЭ��� �����P[Э�P�[�ݭ�������P[Э�P�[�(,����� �e����P�����Э�PЭ��ݬ��~����P[Э�P�[�(,��ЬPݠ��   �ݏ�� ��(          ^� �����P��ݬ��.���(,`��� ������P��ݬ�����(,`��� ������P��(,���Э�PЭ�����Э�PЭ��ѼѼ������Ѽ���Ѽ
���ֽ�ѼѼ
(,���(,���     ^ЬPѰ!+� �L����P��(,���Э�PЬQС����ЬPЭ��        ^� ЬPРPݠ��K����P��� ������P��(,���� ������P��ЬPРP(,������Э�PЭ��Э�PЬQСQС�Э�PРPЭ����ЬPЭ��ЬPЭ��        ^ЬPРPݠ���  �P�P1� � ЬPРPݠ������P��� �Q����P��Э�PЭ�QС����Э�PЭ��Э�PЬQСQС�� �����P��(,���Э�PРPЭ����ЬPЭ��ЬPЭ���P      ^�ݬ������ݏ�� ��%           ^��M�  �,T	 � �   ߬ݬ��3�  ��  �P�%�  ���� � �r         ^Ь[ЬZ�ZH����  �,X	 � �G   ���  �,X	 Y�ZY�ZY�Y�[��͜  ��"  �Yￜ  �Y[�YZ���i� � �           ^Ï,D	   [M��?� $ݏ�� �[�Џ,D	 �p�  ��j�  ��#  !�[Џ,D	 �T�  ��N�  �  ~��L'           ^߬ݬݬ��    �    ^Ь[ЬZЬY��X1� �XP1� ��X�XPe݉�[���   �P[1� ЉW�g����1� ݉�[��"  �P[}݉�[��b  �P[m�YP�Y�`�b�X�]��%��X��X�[�[PtH�P#��P%��P�c   ��P�d   1|��P�l   ��P�o   ��P�s   1o��P�x   ������ �X��X��P#����3��1��k�[P       ^Ь[ЬZЏ�� Y�Z!�ZZ�Z�ݏ�� �[��   �[P6�-�щZ��Y�Y�i�iZX�iXP�PZ�XP�0P��ZP�0P��k�[P         ^Ь[ЬZ�Y�I�ʚ  �I���  Z�Y��Y�Y Q�YQZQ�QP���P�0P��Y�k�[P        ^Ь[ЬZ�Y�I連  �I  Z�Y��YY�YY�Y Q�YQZPʏ����P��� ��Y�k�[P      ^Ь[ЬZ��9m  ���/ ���/ �Z�[ݏ � ��E   ˏ ���[PǏp  PQďp  Q�QPQ�Q���c QX�XYթ�Z�
�[i����Ï�c YP�PO�i[��
Pʏ����P�PZÏ�c YP�P-�Y�Y��� Џ�c Y�YP�YP�PX�ݏH� ����   ^Ь[�X�k�XXP��Q�QPX�ˏ ���XPǏ�  PQď�  Q�QPQ�Q��Џ(� V�V1� �VYЭ�X�W�W��  \�X��  �  X�XXP�PP�YPZ�jݬ�j��X"  �P#�jPOѦ��  ֦ݬ��8   �Pj1�WX�W��fݏ�  ���  �Pf�fV1m�ݏZ� ���      ^Ь[�[��R"  �PZ�Z��" /��   Z��" ��" ��  �P�" ݏu� ��F����Z�[��" ��  �P[�Z�" �Z�" �[P         ^        ^լݏ�� ������ݏ�   ݬݏ�� ���!  ݬ��!  �P��   ݏ�� �ￚ��Џ�� P        ^ݬݬݏ� ������         ^ݬݏ)� ������        ^ݬݏ/� ��������� ݬݏ9� �����        ^ݬ�����լݬݏC� ��t������ 3��y	 ��s	 ݏR� ��R�����_	 PxP~ݏ[� ��9���� ����ݏm� ��%���      ^��P�P�P�Pݬݏs� �酪����Ѭ8Ѭ��Ѭ��ݬݏ�� ��n���ݬݏ�� �����       ^լݏ�� �����2��ݏ�� �����ݏ�� ��u���ݬݏ�� ��e���      ^ݬݏ�� ��K���       ^Ь[ˏ����[P�[P
Џ   P1� �[PU�P1� �P{Џ   Pr�PmЏ   PdЏ�   P[Џ@   PRЏ   PI�PD�P?� P:Џ    P1�P����������������  �����������[ݏ(� ��A���     ^�[�[�K�� �[�     ^Ь[ЬZ���z  *�K�ĕ  ݏ3� ��#  �Z��Zy��ݏ?� ��  �[:�K�� �Z �P�P�P!�[P�PݏC� �ﭗ���[P�@��       ^Ь[x[P�P� �['� �� P� P�P�� P� �� P�PxP�� ��� שּ ���  �� P        ^�[�[�K�� ݏP� ������[�      ^Ь[�Z�k8ݫ<�������PZЫ@[�0�!� ZP� P�PZP
� ZP�PxPZ��@   Z1� ӏ  �� ZP� P�PZP
� ZP�PxPZ� Zkӏ   �� ZP� P�PZP
� ZP�PxPZ� ZEӏ   �!� �4P� P�P�4P� �4P�PxP�4��4Z� ZP� P�PZP
� ZP�PxPZ� Z�ZP       ^��� �P�P�P�Y� ߬ݬ�� ��ݭ�������P�z ��t � � ݏ�� ��Е�����        ^��I Ï � �> ~ݏ � ��@���        ^ЬPѠ
ЬP��	P�P�ݬݬ��6����P��Э�P          ^ݬ������P� Q�QP       ^ЬPݏ�� �� ����P4�P0�P�������������������������������������������       ^ݬ��  �P��լ$Э���խ�����P��P����Q�a`׭��$ά��ѭ�������P��P����Q�a`֭��        ^ݏ�� �龎 ������Ï�  PǏ   PQ�Q����    ��������u� ��  � �  Э�P       ^ЬPcЏ�� Py�  Pp�  Pg�  P^�  PU�  PL��}�  PC��x�  P:��s�  P1��n�  P(��i�  P�P�P   	��������������������1~�        ^��� �Lݏ�� ��PxPP��� P~��R  ���PxPP��� P~��]�����PxPP�(�� ЬP1� �� �.���PxPP��� P~��&�����PxPP�*�� ЬP��PxPP��� (.���PxPP��� P~��������PxPP�*�� ЬP@��PxPP��� $#ݏ������PxPP��� P~�����ЬP�� �ЬP       ^��PxPP��� (?ݏ������PxPP��� P~��Y����)��PxPP��� P~��x
  �`ЬP1���PxPP��� (Ь����PxPP��� �_K��PxPP��� P~ݏ�� �������	��� �
ݏ�� ��PxPP��� P~��M  ЬP1&��PxPP��� �_Ь����PxPP��� *}�+��PxPP��� P~��	  �P��խ��-��PxPP��� P~��	  �P��խ�Э�P��
Э�P��(1� ݏ������PxPP��� P~��!���ЬP��PxPP��� *Ь�1j���PxPP��� �L.���PxPP��� P~��������PxPP�&�� ЬP&��PxPP��� �LЬ��ݏ�� ���         ^��� �
ЬP1� ��� �ЬP1� ��
ЬP1� ��ЬP1� �� �
ЬP1� �� �ЬP1� �-��PxPP��� P~��X  �P#�+��PxPP��� P~��;  �PЬPL�-��PxPP��� P~��  �P#�+��PxPP��� P~���  �PЬP��  �
ЬP       ^ѼЬPѰ2�P1� �P1� мPTݏ � ��Y���ЬPݠ������PЬPݠ������P�P�P1� ЬPݠ�����v�Pr�Pm�P2������������������������������������������������������������������������������������������������������1?�     ^� �����P��мP1_ЬPݠ<�������P��ЬPݠ@�������P��Э�PЭ��Э�PЭ��1ЬPݠ<������P��ЬPݠ@������P��Э�PЬQ2�:�(Э�PЭ��Э�PЭ��1�ЬPݠ<��X����P��ЬPݠ@��F����P��Э�PЬQС4�$Э�PЭ��Э�PЭ��1�ЬPݠ<������P��Э�PЬQС4�Э�PЬQС8� Э�PЭ��1XЬPݠ<�������P��Э�PЭ��Э�PЬQС@�Э�PЬQС4�$1 Э�PЬQС4�Э�PЬQС<�Э�PЬQС@�1� �P�v   ��� ��� ��������^�����^�����^���������� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� ��������������������� � ��� ^�� � � � ^������ � � � � � � � � � � � � � ��� � � ������ ^���^�� � � ^�� ^���^�^�� ^�����������мP1rݏ
� �� ������1W���1P���1I���1B���1;���14���1-���1&�	��1�
��1���1���1
���1���1����1����1����1����1����1����1����1����1����1����1����1����1����1����1����1����1����1�� ��1~�!��1w�"��1p�#��1i�$��1b�%��1[�&��1T�'��1M�(��1F�)��1?�*��18�+��11�,��1*�-��1#�.��1�/��1�0��1�1��1�2��1 �3��1� �P�v   ��������&��������
��������������������������������������������������������������������������������������B���;���������������4�-�����I�������������^�����������������������������������������W���P�������e�������s���l���z�����������������1��ЬPРP1� ݏ� �憎��Э�P��1Э�P��1Э�P��1Э�P��1� Э�P��1� Э�P��1� Э�P��1� Э�P��1� Э�PԠ1� Э�P�	�1� Э�P�
�1� Э�P��1� Э�P��1� �P��   �B�P��P1n��P1N�1>��P�16��P ��P�1'��P�@   13�1��P�   1q�,�P�   1B��P�   1J�1���P�   1f�1���P�    1b�1��1��        ^мPW�P1� ЬPݠ�������PЬPݠ�������P�P�P1� ЬPݠ������P{ݏ3� �����l�P2�������������������������������������������������������������������������������������������������������       ^ݬݬ���            ^ݬݬ��            ^ݏJ� ��^��� ��V� �M�    �     P      �ЬX��X�SЬR�U��T� T��T�T�+T�-T�S��T|P�T04�T9/�Q����yPVyPP�VP�WQ�0T�TP� Q�U�S�U��TǑT.�S��V�T�e�T�E[��T�T+�T-�S��T�T0�T9�V������FfV>F��V��S�VV�VU�U�����Џ����U�U�d   Џd   U�X�R�Rh}PP1� �R�U#�Q����	y��PP�R�yPV�VP�WQ�R�U�=;�QyPP�RyPP�R�Q��QV�W{VQW�PV� W{
VPV�PP�V�P�R� U��Qy��PP�RyPP���PPnPVnQPd�~���P`VP� SrPP�RpP~��     � ^Ĭ�ݬ��L  �P[ݬ� �[��=  �[P      � ^ݬ���    ��h  �P   � ^� �   ݬ������  �^Ь[�  �  ��C  ��  �����������.Џ����P1� ЫZi�[��� 9�� ���� ����� ���א����X�X߭���~��~  �PY�kVݏ   ��^  �PZ�Z�������Y�YX �Z�Y�YX�Z��Y�Z��~��3  �PYЏ�  k����Z��XY� �1L�ЬP    � ^Ь[2�Pʏ����P�PHЫZB�Z�Y;�Z���� ��PЏ   P�Pk�Y�Z��~��  �PY� �Џ����P�P    � ^�渚  [�����	�[��t����[�[��  �    � ^Ь[Џ����Z���A��<�[��>����PZ��~������PЏ����Z��
ݫ���  ��� �ԫ�����k�ZP      ^ЬP���� �ݬ���  ݬ߬ݬ���  �P[ЬP�� �QѠQݬ������ ݬ��  ЬP��	Џ����P�[P  � ^Ь[ЬZ��+�P�P�PX�k�w+ݏ�  ݬ��
  �PY�X1� �Y��Y��"����{�k�aj�X�~�~ݬ��  �PY<��_� 3ݏ�  ݬ��d
  �PY�X�Y�Y�������ݬ��L  �PY�Y'�� �Y���   �X�~�~ݬ��!  �PY�Z��I����Y�P&�j�Y��X���k�r�����ZP     �^߭�ݏt  ݬ��  �P
��� �P�P   p�P�PR��R�R�   
�RP|Pp�ȋ  P��rPP�"�\�      ��X	      � ^���~��  �PZ�Z  J�Z8�ZP�P�PZP�PP�PP�@�t Y�i['�kP�[P�P�ZP�[�ki�[P� ��  ��W�  �Z��        � ^Ь[��1�  Z�X�j3�Z�$�  �ij�jY�i��[[P�PP�ZP�YP�[[P�PP�ZP�PZ1� �ZY�jZ�ZY��X�X	��ۊ  Z�� ���  �PZݏ   ��   [~��  x
PX�XXP�PP�ZP�PZxX~��  �PY�Y�����&�[XP�P�PX�[XP�P�� �  �P19��P1x � �  xX~�Y��7  1��[[P�PP�P�F�  �Y�?�  ��7�  �& �j�+�  ��$�  j�Z��  	�Y��  ���  ����  Y�Y���  ��ZP    � ^Ь[]�[�kP�[P�PY�Y�؉  ;�Y6�YP�P�PYP�PP�PP�@� X�hZ�jP�ZP�P�YP	�Z��[h�[~��       � ^Ь[�[�[�q�  �[�f�  �[�]�  �k� �^��} [ԭ��Z�Z�����֭��jk�kZ��[�[�8X	 �Э�P   �^ЬZ�ݬ��  �PP�PP�ZP�P��Э�j�Z���  W���  [��ۈ  YЭ��ވ  �[P�ZP�ZP�ZP�Pk���P�YP�YP�YP�P������    ����  ���^Ь[ݬ������1� ��	�[�������[��P�P�����~��_  �PW�W~������PX�X[�XPN�W���W���[Z�XYЊ�Э�P׭��P��X[��WWP�PP�XP�P[��WWP�PP�XP�[P�P��� @h�     � ^  @ ЬV#}�S�TQя��  V(���ac��  V�(VacЬP� ЬV'}�S�TWя��  V, lW���c��  V�, lWVcЬP  �^ԭ�Э�P�@�� Ь@��� �P	�!����P      ���         ^��  �� ���  ��^  ��  ߬ݬ��I  �P[�� �P��y  P��h  ��5���� ��Y  ��  ��W  	Џ����P�[P     �^Ь[ЬZԭ�լ05Ь���jЪP֪�`P	�Z��  �PY�Y�׭��֭�ѭ���Э�P   �^Ь[ЬZԭ�լ16ЬY�j��PЪQ֪�Pa�Z��~������Y���
֭�ѭ���Э�P   ��       �������  �~��\S�^\��  ���  P����    ��g  Ь�υ  �P � ^Ь[�  �  ��S��������ի��
ݫ�������� �Ь���Ы��k   ЬPЭ`Э��P  ЬP�PЬQ�aP���P����Q�
���Q��a�(Џ�U ����7   ��   ��^�С��ݏ[V ���:   longjmp botch
    �0�d      �^��B ��Ь��Џ�  ��߭�߬ݬ���  �P[׭��PЭ�Q֭��Pa߭�� �������[P �Џ��  X}�V�VQ: Xa��QS: Xg(Xgc�QW������WQ�Q(Qgc�VP     }�R: ���b:S���b�QR������RQT�T:STb�QP   }�S�ST�P: ���d)���dc�QT������TQ�Q)Qdc�acP�PP  � }�V�VS: ���g(���gc�QW������WQ�Q(Qgc�VP     ЬR�RQ: ���a��RQP  �ЬUC}�S�TV�URЏ��  Y�YUX�YU: Uf�VQU�X�YRW�YR,Uf Rc�WR	�XU��U�ЬP � ^Ь[��Z�Y�kZ�[Y����YP      �ЬQ�Pa  �#   ЬPЬR�R�Q{RPPR�PR�P�P   ЬPЬR�R�Q{RPRP�P�PR�RP   ��<        �^� ��$Э�P�@�� �@�� ���@�� � ��׭�խ��   �P��� �P   ������    	
 !"#$ &'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������T7��R�B�����d�ݭ��R��z����P��� ֭�������S}��T�T��P���R�P�T��S�C�����R�Q�S��T�P�}T���P���R�P��P�Q�R��� Э�P��� �^Ь[Ь��Ь\ԭ�<���P�[Q}��T�QUR�PR�RP0r��Q[�Rܕ���^U|Y|V��P�P �X�� � �� � � � � � ��� ��� ����������� � � � � � � � � � �� � � � � � � � � � � � � � � y� � � � � � � � � � � � � ��$���� � � ��� � � � � � � y� � �P�1��1�ȏ@   Z� P11��XP�Z�PЌR: Pb�QU�RQ1'0123456789abcdef0123456789ABCDEF�R�S������W�R�S������W�Z������W�SV�Q�UЌP�RSPQ�Ag�� VR��|V�e;0��Z1} լ�1u �S��xP�Z��XP�Pq�W�0qYʏ�   Z�lP�P
n4
n� 
�
n� ��   
n� ��
n�W8
n������; ��W�Z�+q�Z� q�W�Z�X�QUV�WV�VX&�WQ�Q�H� R�]R�RX(VaHa, a0X� �W�Q�VSU�QUX�XYP �Z�ZR�WP	�PX�PY0)��XYP7�XY�XP0��R�P��R}��T�T0���R�֭�}T����YP1b�1]��0R� R�PY�Q�PW�P^, `RWn�WP�^Q0���W^ЎQЌP�P��^Q1i�ȏ�   Z1L�� Z1F��Z1@��Z1:�� Z�Z�Z�Z�IiY>I��Y	�HhX>H��X�Z1��X�Z�Z1��ZЌY��Z�YY�ЌX��XX��Z�X0����XW�WV�W�W�W�WP�PnW�#� V�WP֭��W�P�H��� W�x��WP���@���Q�WV��S�����0��0S��, a��Vc�c8Va�0��VUQ�nS�W���-��WЭ�P�0��PV�VP�PV�P��(PacЭ�P, a0Pc�XP�Z�	Z�.�έ�P�PX�XP�PX, a0Pc�XP�PV�VP�PX(Pac�XP�@� R�]R�RP�PX�PX, a0Pc�SU�DeB+� �X�Z�X0� �XW�W�W�WP�PnW�֭��WP�P�=��� W�x��WP���@��Z=��Q&�QV���P�Pn8n����e�VQ�Z1,�� ��1%��WV�XЭ������1�����P0�P�PX(�WV�PX��Q0���Z�	Z�u0��e.�U�Z�1����Q0���Z��Z�X�X�X�Z1.�1+����p�U1� rUU����UR���R�;R��� R���RƏ�   R0� qPU�R�R���RR�R
d��   U�R�	R�\   tPTUPU�P	��	� �t�    UPU�P��XW�����юn���W�W	qU �� ������P����   pP�T~�M   S�R�RR�R �TRdcP�S�T��RgPP�R������Q�RR�(RS�S�A   �����Q�B�b   T B      �C      G @    �M �    [��  �u��+��pPB<�   �Vvӈ�b��2>H�QS'���I[��������#,;
�                         ��:��ܒ� �X��  � ^Ь[�����
Џ����P1� ���ݏ   �������P���ի��ߘ�P�@�� ����[��� ���q  ���q  ��������~Џ   ~ݫ��~��(����PkЫ��k!�k���������
��� ��k1Q�ЫP֫�`P     �6����                                                                                                                                                                                                                                                                                                                                                                                                                                                               @(#) cgram.y:	2.1 83/08/02      ��   ��    2  9  ��  �� 8 P 9 P �� �� 3 D ��B �� : M ��O �� : N ��S ��" 4 + ��) ��$ 4 # ��! ��8 5 / 9 / ��  � � F  " 
  N ^ e �  c � Z X Y  � Q  b O � � P    7 ] ` � g :   7  S R 2 A 6� � � L � � � � � � � � T d U ,m �  o � � %� 	 � k   � &   � c � � � � � � � � b K j � � \ h & % 4 ` 8 � p  � f � q � � � � � � � � � � � � � � � � � d r � n  � � � � � � � � � � � � W Z X Y ( D J � ) � * , ( � 8 � ) � 0 � 0 � 1 � 1 � � � S R � @ � � 0 C � c 1 � � � _ � # T b U ! :� � � �   
  � � � � ) �  � � � I   m   H ? � � � � +* d , 	
  _  
  �  G W Z X Y Q  !O a � P # � � 3 
 5   &'  y S R  *� Z X Y � Q i  O 0u P T  U #� 5; 4$ #" B ;9S R � + - 8� � � 1� � � � � � � � T 2U a m _ l v � w � � y  < { / E | . } � � � ~  � s z u x v [ w 6 9 y � v { w � | y } > � = ~  � s z u x ' � t s � u x   � V  v  w   y   { 3� | � } t � � ~  � s z u x v � w �  y             v   w     y     { /u |   } t � � ~  � s z u x                         v   w     y     { .  |   } t � � ~  � s z u x   v   w     y               v   w     y   -{ u x | t } � � (~  � s z u x v   w     y �   {     |   }   �   ~  � s z u x   v t w �   y     {     |   }   �   ~  � s z u x   t $�                         v   w     y     { t | � }   �   ~  � s z u x v   w     y     {     |   }   � � ~  � s z u x     t �               v   w   v y w   { y   | { } t � � ~  � s z u x s z u x                 v   w     y     { �   |   } t � � ~  � s z u x v   w     y     {     |   }   �   ~  � s z u x     t   � W Z X Y     Q     O     P W Z X Y     Q     O �   P     S R                       S R       T   U     W Z X Y   � Q   T O U   P W Z X Y   � Q     O     P     S R                       S R       T   U     W Z X Y   � Q   T O U   P W Z X Y   � Q     O     P     S R                       S R       T   U     W Z X Y   � Q   T O U   P W Z X Y   � Q     O     P     S R                       S R       T   U     W Z X Y   � Q   T O U   P   W Z X Y �   Q     O     P   S R   v   w   v y w   { y   S R }  T  U   � s z u x s z u x   T  U W Z X Y     Q     O     P W Z X Y     Q     O     P     S R                       S R       T   U   M W Z X Y     Q   T O U � P W Z X Y     Q     O     P     S R     v   w     y     { S R |   } T � U ~    s z u x     v T w �   y     {     |   }       ~     s z u x v   w     y     {     |   }             s z u x ������4  �� � �� ��� 8� 5��. q �� � �y ���� �� � � �3�����  y q � i   � � f ����+ �S 7 ��� �� ��Q ,��9 �����O ��r ,,,,,9�� ���� � 6 �w ��� �� � 3��q � �����1�,,��aT.,!��,,,,, �����,%�r r r r r r �� �� �8 ����������* �� ����,,,�,�,q�,�,�,zbm��� � R�� ,�_ � � ,�S ��  ��������,��� �,� r < �^ _ ��� ��U& �  � �    � $��� � �� � ,	H�-�; � ���� �� � ,���� ���,,������ �,�  ��������,����j, �������,�  �  �. �������     �H ��  �	 )� ��� ��~"   z v t
 $ sq' fdba( _^  \WVQGC@;               ! ! # # #        $          % % ' '     ( ( * *   +                  ,  .  	 - - -  0  1 1 / / / / / 2 2 3 3 & & ) ) 4  5 " " " " " 6 7 " " 8 9 " " " " " " " " " " " : : :     ;      
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
                                                                                                                                                                                                                                          ������� ; ��������" ! ������# ��1 9 9 ������ 2 ������  ����! 4  4  9 8 ��2 6 ������������2 6 : 2 ��! ���������� ������3 7 ����3 3 ��  3 3 7 ����4 ��     0 2 ��    ��9 ������    2 ��8 : ����������4 7 ��3 8 7  8              : ��������4  6   2 ������������2 ������3 ����2 5 ��8  ��5 ������9 �� ������: ��: ��: ��: ��: ����: ��: ��: ������������8 ���� ��3 3 ��2  8 3 ����9 �������������������� 5 ����7  3 ��6 3 ��������9 ����5 ��; ������+ ��- ��) * $ % 9  ��& , (  / . ��5 ��7 ��3 9 9 9 ��������2 ��9 9 9 �� 9 5 ��2 2  �� 7 7 2 ' 2 + ����9 9 ���� 3 ��2 9 3 3 3 ������3 ����9 9 ����3 �� ��                *   "     ��J     ����  ��;      ��  �� K    | 7 =           |   F   Z , ��X $ &   	   > ?     < A   G I E 8 9   Q   �                 � � � �   [ . 0 3 | 6   ;     Y | L P 
    ^ @ } C   :                                 X T V   \ �     � � � � � � �       � �   � � ( - 1 | 5   % '     H � � �   �   �   �   �   � �   �   �   � �   � �   Y X   �     � � � �   �   4      � � � � � � � �   R U   �   � � | �   � � 2     ]     a     d               q       x   �     � W   �   �  _ ` b c      k l m n     r s t     u   w � �   z       ~ o p     v �     h y { e          f g i      j         P� U� \� a� f�     h�         j�         l�         n�     p�     r� t� v� y� |� �� �� �� �� �� �� �� �� �� �� Ê ʊ ϊ Ҋ ׊ ފ � � � �� �� � � � � � � � � � � !� #� %�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             )� *� K� L� M� N� b� ~� � �� �� �� �� �� �� �� �� �� �� �� �� ΋ ϋ Ћ � � � �  � !� "� #� $� %� C� D� \� ]� ^� _� `� l� m� n� o� �� �� �� �� ƌ ǌ � � � �� �� �� (� )� *� +� E� F� n� o� p� |� �� �� �� �� �� �� �� �� �� �� �� ٍ ڍ � �� � $� :� n� �� �� �� �� �� ��  Î Ď Ŏ Ǝ ǎ Ȏ � � �� � � � � � � :� ;� <� =� >� ?� _� `� q� ~� �� ɏ � � ;� L� n� �� �� �� ̐ ݐ � �� �� �� �� � � � I� c� d� e� f� g� h� i� j� �� ё �� �� �� � � � � � � � � � � � (� )� *� +� ,� -� .� A� B� Q� R� a� b� w� x� �� �� �� �� �� �� �� �� �� �� ޒ ߒ �� �� �� �� !� "� .� K� L� M� N� O� d� e� �� �� �� �� � �� �� �� �� �� �� �� �� � � � � � 4� 5� 6� 7� 8� I� J� K� L� M� e� f� g� �� �� �� � 	� 
� :� e� �� �� �� � � � 4� S� j� k� �� �� �� �� �� �� ϖ Ж � �� �� �� �� �� �� � O� P� Q� R� S� T� q� �� �� �� �� �� × ė � � � � � � +� [� �� �� �� �� �� �� �� �� Ә � � � � � �  � E� u� �� �� �� �� �� ϙ ��     ����        bad bdty dimension table overflow whiles, fors, etc. too deeply nested non-constant case expression case not in switch switch table overflow duplicate default in switch default not inside switch switch table overflow duplicate case in switch, %d char %d in %s %s in %s yacc stack overflow lex EOF
 lex %s
 lex (%c)
 lex EOF
 lex %s
 syntax error
%s saw %s
 saw `%c'
 saw EOF
 saw char 0%o
 error recovery pops state %d, uncovers %d
 error recovery discards  %s
 `%c'
 EOF
 char 0%o
 reduce %d in:
	 function level error $%dFAKE union member must be named field outside of structure illegal field size field outside of structure zero or negative subscript arg list in declaration function declaration in bad context arg list in declaration nesting too deep loop not entered at top bad while loop code gen value bad while loop code gen. value loop not entered at top bad for loop code gen. value bad for loop code gen. value illegal break illegal continue statement not reached void function %s cannot return value loop not entered at top precedence confusion possible: parenthesize! old-fashioned assignment operator & before array or function: ignored structure reference must be addressable undeclared initializer name %s  NAME STRING ICON FCON + - * & | ^ ? : && || ASGOP RELOP EQUOP DIVOP SHIFTOP INCROP UNARYOP STROP TYPE CLASS STRUCT RETURN GOTO IF ELSE SWITCH BREAK CONTINUE WHILE DO FOR DEFAULT CASE SIZEOF ENUM ( ) { } [ ] , ; = ASM  expected an external definition
    semicolon required
 expected one of NAME * ( ;
        { expected in struct decl
  { expected in enum decl
    expected , or ;
   expected one of NAME * (
 expected one of NAME * (
   expected = in intializer
      expected TYPE STRUCT or ENUM
  an enum must be a NAME
     ) required
    expected ( ) or [
 expected ( ) or [
 expected a NAME in list
 ) required
 ) required
  { or expression required in intialization
      type_declaration expected one of NAME * : ( } ;
    expected one of NAME * (
  function_body needs a declaration or {
   ] required
 need constant expression
   expect ) or ,
      ] needed
  expecte expr or { in initializer
  term :  *.term 
 term :  &.term 
 term :  -.term 
 term :  UNARYOP.term 
 term :  INCROP.term 
 term :  SIZEOF.term 
term :  SIZEOF.( cast_type ) 
 term :  (.cast_type ) term 
term :  (.e ) 
 expected ) or expression
     } needed
       expected one of NAME * (
  expected one of NAME * (
 enum_dcl must end with }
      expected one of NAME * : ( ;
      name_list :  name_list ,.NAME 
  e :  e RELOP.e 
 e :  e ,.e 
 e :  e DIVOP.e 
e :  e DIVOP.ASSIGN e 
 e :  e +.e 
e :  e PLUS.ASSIGN e 
 e :  e -.e 
e :  e MINUS.ASSIGN e 
 e :  e SHIFTOP.e 
e :  e SHIFTOP.ASSIGN e 
 e :  e *.e 
e :  e MUL.ASSIGN e 
 e :  e EQUOP.e 
 e :  e &.e 
e :  e AND.ASSIGN e 
 e :  e |.e 
e :  e OR.ASSIGN e 
 e :  e ^.e 
e :  e ER.ASSIGN e 
 e :  e &&.e 
 e :  e ||.e 
 e :  e ?.e : e 
 e :  e ASOP.e 
 e :  e =.e 
    initializer needs expr or {
   term :  term [.e ] 
term :  term [.e : e ] 
 term :  term STROP.NAME 
        term :  (.cast_type ) term 
term :  SIZEOF (.cast_type ) 
term :  (.e ) 
 term :  ( cast_type.) term 
 expected operator or ) after expression
   expected , or )
           expected , or ;
       e :  e DIVOP =.e 
  e :  e + =.e 
  e :  e - =.e 
  e :  e SHIFTOP =.e 
  e :  e * =.e 
   e :  e & =.e 
  e :  e | =.e 
  e :  e ^ =.e 
   operator expected after expression
   init list must end with }
   operator expected after expression
  ) required
 term :  ( cast_type ).term 
     elist :  elist ,.e 
  expected one of NAME * : (
   expected one of NAME * ( ;
 stmt_list :  stmt_list.statement 
compoundstmt :  begin dcl_stat_list stmt_list.} 
         e :  e ? e :.e 
   } expected
  term :  term [ e :.e ] 
     expected ) or [
     expected one of , or ;
   ; or operator expected after expression
 ; reuired
  statement :  ifprefix.statement 
ifelprefix :  ifprefix.statement ELSE 
 statement :  ifelprefix.statement 
  statement :  doprefix.statement WHILE ( e ) ; 
 statement :  FOR.( e ; e ; e ) statement 
 statement :  switchpart.statement 
 statement :  BREAK.; 
 statement :  CONTINUE.; 
 statement :  RETURN.; 
statement :  RETURN.e ; 
 statement :  GOTO.NAME ; 
  statement :  error.; 
statement :  error.} 
 statement :  label.statement 
 ifprefix :  IF.( e ) 
  switchpart :  SWITCH.( e ) 
  label :  CASE.e : 
 label :  DEFAULT.: 
   expected an operator or ]
  null_decl :  null_decl [ con_e.] 
       statement :  WHILE .( e ) statement 
 statement :  doprefix statement.WHILE ( e ) ; 
      expected a ; or an operator
 statement :  GOTO NAME.; 
    ifprefix :  IF (.e ) 
 switchpart :  SWITCH (.e ) 
  expected a : or an operator
    null_decl :  ( null_decl ) (.) 
  statement :  WHILE (.e ) statement 
 statement :  doprefix statement WHILE.( e ) ; 
 statement :  FOR ( e.; e ; e ) statement 
    expected ) or operator
 expected ) or operator
   expected ) or operator
 statement :  doprefix statement WHILE (.e ) ; 
     expected ) or operator
  statement :  WHILE ( e ).statement 
 statement :  doprefix statement WHILE ( e ).; 
 statement :  FOR ( e ; e.; e ) statement 
     statement :  FOR ( e ; e ; e.) statement 
 statement :  FOR ( e ; e ; e ).statement 
                           ����p� t� z� � �� �� �� �� �� �� �� �� �� �� Ś ͚ ՚ ۚ ߚ � FIELD[%d]   SNULL AUTO EXTERN STATIC REGISTER EXTDEF LABEL ULABEL MOS PARAM STNAME MOU UNAME TYPEDEF FORTRAN ENAME MOE UFORTRAN USTATIC                     t2	 t2	 $       _      0             
      "      '      `      (  2   )  3   {  4   }  5   [  6   ]  7   *    ?     :     + 	   - 
   /   < %   > &    |    ^    !   L ~   M ,  8 8 ;  9   .    D <   S >   U =  : : ��     �        �       !�    )   '�    /   ,�        1�    *   :�    .   B�    ,   E�        L�    '   Q�    1   V�       ]�        c�    -   g�       o�    %   t�    &   w�        {�        ��       ��    $   ��        ��    0   ��       ��        ��    (   ��       ��        ��        ɠ        Π    +               bad option: X%c ccom: can't open %s
 w ccom: can't open %s
 %s -- line %d %s
 # %s %s # abcdefghijklmnopqrstuvwxyzABCDEFGHIJKLMNOPQRSTUVWXYZ_ 0123456789 0123456789abcdefABCDEF  	 01234567 abcdefghijklmnopqrstuvwxyzABCDEFGHIJKLMNOPQRSTUVWXYZ 123456789 	 lxstr() unexpected EOF newline in string or char constant non-null byte ignored in string initializer empty character constant too many characters in character constant lxcom() unexpected EOF illegal character: %03o (octal) illegal hex constant yylex error, character %03o (octal) out of switch in yylex asm > %d chars bad asm construction bad AR_?? action %s
%s
%s
 #ASM #ASMEND    asm auto break case char continue default do double else enum extern float for fortran goto if int long register return short sizeof static struct switch typedef union unsigned void while             defid call tyreduce defid( %s (%d),  , %s, (%d,%d) ), level %d
 	modified to  , %s
 	previous def'n:  , %s, (%d,%d) ), level %d
 declared argument %s is missing 	previous class: %s
 redeclaration of: %s from line %d redeclaration of %s from some line %d 	new entry made
 void type for %s too many nesting levels (%d>=%d) 	dimoff, sizoff, offset: %d, %d, %d
 too many arguments (%d>=%d) parameter stack overflow (%d>=%d) bcsave error parameter reset error switch error dclargs()
 	%s (%d)  
 %s$%d.%d dclstruct( %szindex = %d
 ?? gummy structure member structure member has size 0: %s zero sized structure 	dimtab[%d,%d,%d,%d] = %d,%d,%d,%d
 	member %s(%d)
 redeclaration of formal parameter, %s compiler takes alignment of function illegal use of function pointer using a void value unknown size too many initializers (%d>%d) inoff error beginit(), curid = %d
 instk((%d, %o,%d,%d, %d)
 no automatic aggregate initialization insane structure member list endinit(), inoff = %d
 too many initializers (%d>%d) empty array declaration %d initializers for a scalar cannot initialize extern or union } expected doinit(%o)
 initialization by non-constant illegal { irbrace(): paramno = %d on entry
 local variables fill memory structure larger than address space local variables fill memory illegal field type field too big (%d>%d) zero size field structure fills memory structure overflows memory nidcl error illegal type combination tymerge: arg 1 array of functions is illegal function returns array or function a function is declared as an argument function illegal in structure or union parameter declared with weird storage classs function has illegal storage class field not in structure illegal class illegal class illegal class register declaration outside a fncn auto outside function illegal class fortran declaration must apply to function fortran function has wrong type illegal class: %d Symbol table full 	nonunique entry for %s from %d to %d
 removing %s = stab[ %d], flags %o level %d
 %s undefined symbol table full %s redefinition hides earlier one 	%d hidden in %d
 unhide uncovered %d from %d
 unhide fails                        9� ?� D� I� O� S� X� ^� e� k� s� z� �� �� �� �� �� �� 
       syntax error: colon in subscript buildtree( %s, %d, %d )
 constant argument to NOT constant in conditional context struct/union in conditional illegal lhs of assignment operator %s undefined %s not struct/union member member %s==%s?
 %s not in this struct/union nonunique name (%s) demands struct/union or struct/union pointer %s needs reference to struct/union undefined structure or union %s not in this struct/union illegal indirection can't take address of cast unacceptable operand of & assignment of different structures type clash in ?: call of non-function call of non-function other code %d chkstr( %s(%d), %d )
 undefined struct/union using %s gummy structure illegal member use: perhaps %s.%s? division by 0 division by 0 division by 0 illegal shift enumeration type clash, operator %s pointer/integer structure pointer array size pointer illegal %s combination, op %s undefined bit field type pointer required structure appears where arithmetic type required union appears where arithmetic type required bad bigsize: 0%o cbigger trying to cast to a struct, void or union illegal oconvert: %d illegal pointer subtraction incompatible types in ?: void type illegal in expression tymatch(%o): %o '%s' %o => %o
 integer constant expected constant too big for cross-compiler no structure casts operands of %s have incompatible types sizeof returns 0 
++++++++
 T ---------
 R 	      %s=%d) %s,  lval=%ld , rval=%d,  type= , dim=%d, siz=%d
 L undef farg char short int long float double strty unionty enumty moety uchar ushort unsigned ulong ? ? PTR  FTN  ARY  %s statement not reached L%d L%d     P Q T U R S X Y V W tydown(%d) called with:
 tydown:
 tydown(%d), after doptim(R):
 tydown(%d), after doptim(L):
 sconvert(%d) called:
 sconvert doptim called on:
 doptim works on:
 optim did
 optim did
 & error optim did
 optim replaces op1 (%d) by:
                              �  �                  giving up
 internal error floating point error 	casel	r0,$%ld,$%ld
 L%d:
 	.word	L%d-L%d
 	cmpl	r0,$%ld
	jeql	L%d
 	jgtr	L%d
 	.space	%d
 incode: field > long 	.long	0x%x,0x%x	# %.20e
 	.long	0x%x	# %.20e
 	.set	L.R%d,0x%x
 	.set	L.SO%d,0x%x
 	.word	L.R%d
 	subl2	$L.SO%d,sp
 	movab	L%d,r0
 	jsb 	mcount
 	.data
 	.align	2
 L%d:	.long	0
 	.text
 	.data
	.comm _proFptr,4
	.text
 	tstl locprof+4
	bneq L%da
 	movl _proFptr,locprof+4
	moval locprof,_proFptr
 #entry %d
 L%da:	incl locprof+%d
 	.globl	%s
 %s:
 	.lcomm	L%d,%d
 	.lcomm	L%d,%ld
 	.lcomm	%s,%ld
 	.comm	%s,%ld
 Non-static/external in common e2print called t2print called             Q   P   U   T   S   R   Y   X   W   V   ����force bad option: %c genbr genbr1 rcomma    E  vaxpcc2 	.stabs	"%s",0x%x,0,%d,%d
  	.stabs	"%s",0x%x,0,%d,%s
  	.stabn	0x%x,0,%d,%d
   	.stabn	0x%x,0,%d,%s
   	.stabd	0x%x,0,%d
  d   L%d %s: unexpected stab class %d: %s, type = 0x%04x
 %s: 	.data
locprof:	.long %d
 	.long 0
	.long L%db
 	.space %d
 L%db:	.byte  0x%x, 0
 	.text
 %s:          ""                                                                                                  `@                                                                                                                                                                                                                                             x�    NAME          STRING     ^   REG        _   TEMP       t   AUTO       u   PARAM         ICON          FCON       `   CCODES     
   U-            STAR          U&         H   UCALL     K   UFCALL    L   !          M   ~          q   INIT       h   CONV          +       h     +=      i!     -       (  	   -=      )!     *       	     *=      	)     &       h      &=      i      ?             :             &&            ||         8   ,          ;   ,OP        a   FREE!?!    :   =       	   <   /       �  =   /=      �!  >   %       �   ?   %=      �   @   <<        A   <<=     	0  B   >>        C   >>=     	0     |       h      |=      i      ^       h      ^=      i   N   ++      	   O   --      	   E   ->         F   CALL      I   FCALL     P   ==         Q   !=         R   <=         S   <          T   >          U   >          Y   UGT        X   UGE        W   ULT        V   ULE        ]   A>>        !   TYPE       6   [          m   CBRANCH    l   GENLAB     p   GENUBR     n   GENBR      o   CMP        g   FLD        i   P*         j   P/         $   RETURN  	   r   CAST    	   %   GOTO       b   STASG      c   STARG      d   STCALL    f   USTCALL   v   RNODE      w   SNODE      x   QNODE      �   MANY       s   ARG        y   UOP0    @  z   UOP1    @  {   UOP2    @  |   UOP3    @  }   UOP4    @  ~   UOP5    @     UOP6    @  �   UOP7    @  �   UOP8    @  �   UOP9    @  ����            %s:%d: 
 too many errors cannot recover from earlier errors: goodbye!
 compiler error:  
 warning:  
 out of tree space; simplify expression wasted space: %d nodes out of temporary string space out of memory [tstr()]           ��    �  ��    �  ��    �  ��       �� �  �  �� ]   �  �� :   �  �� F   F   �� I   F   �� H   �  �� K      � m   �  � 8   �  � o   �  !�    �  &� ;   �  ,� M      2� h      8� �  �  =� O   �  B� <   �  G� =   �  K� �  �  R� �   �   X�    �  _�    �  b�       h� g   g   m� s      q� a   a   x� n   n   }� l   l   �� p   l   �� %   %   ��       �� N   �  �� q      �� �   %   �� �  �  �� @   �  �� A   �  �� �  �  ��    �  �� 	   �  �� 
      �� >   �  �� ?   �  ��    �  ��    �  ��       �� L      ��    �  ��    �   �    �  �    �  �    �  � �   �   �    �   � ^   ^   &� P   �  *� Q   �  .� U   �  2� T   �  6� S   �  :� R   �  >� Y   �  B� X   �  G� W   �  L� V   �  Q� $   $   V� &   �  ]� v   �  i� x   �  o� w   �  u� B   �  {� C   �  ~�       ��       �� c   c   �� b   b   �� E   b   �� d   d   �� f   �  �� �   �   �� �   �   �� �   �   �� �   �   �� _   _   �� t   t   �� u   t   ��                 #tree  ??? (unk op %d ???)  (%s %d???)  )  )  )  %d)   %d %d)   %d %d  )  %d  )  )  %g)   %s L%d  )   L%d  )   L%d  )  %s+%d)  %s)  %d)  %d)  %s+%d)  %s)  %s)  L%d)  %s %d)  %s)  %s   %d L%d)   L%d)   %d %d)   %d %d  )   %d  )   %d %d  )  %d  )  %d)  prtype(#%x)
 C UC S US I U L UL F D St P %s  #treeend
   ??? and andand asgand unaryand arg ars assign call fortcall unarycall unaryfortcall cbranch  cm  cmp  colon comop compl conv copy decr div asgdiv entry epilog er asger fcon fld funarg free genbr genlab genubr goto icon incr init labelpt locctr ls asgls lxinfo minus asgminus unaryminus mod asgmod mul asgmul name not or asgor oror  plus asgplus prolog quest reg eql neq gtr geq lss leq gtru gequ lssu lequ return unaryreturn rnode qnode snode rs asgrs star star starg stasg stref stcall unarystcall swbeg swcase swdef swend temp vauto vparam   #	reg	%d
 expression too complicated #	incl	locprof+%d
 codegen failed at top level #%d  
 #	weird??? %d
 #	bit%c	%s,%s
 $%d #	mcom%c	%s,%s
 #	bic%c2	%s,%s
 #	bic%c2	%s,%s
 #	bic%c3	%s,%s,%s
 %d arguments is too many #	calls	$%d,%s
 ) #	push%c	%s
 #	clr%c	%s
 #	cvt%c%c	%s,%s
 #	cvt%cl	%s,-(sp)
 #	mov%c	%s,%s
 #	cmp%c	%s,%s
 #	mcom%c	%s,%s
 movz cvt #	mov%c	%s,%s
 #	%s%c%c	%s,%s
 #	mov%c	%s,%s
 sub no float ++/-- #	mov%c	%s,%s
 inc dec #	%s%c	%s
 #	%s%c2	%s,%s
 (%s) *%s weird asaddr in incrop inc dec #	%s%c	%s
 #	%s%c2	%s,%s
 div udiv xor #	%s%c3	%s,%s,%s
 #	mov%c	%s,%s
 #	cvt%c%c	%s,%s
 #	inc%c	%s
 #	dec%c	%s
 #	%s%c2	%s,%s
 #	push%c	%s
 #	%s%c2	%s,%s
 #	%s%c3	%s,%s,%s
 ) #	mov%c	%s,%s
 #	ext%sv	$%d,$%d,%s,%s
 z  #	%s	 #	tst%c	%s
	%s	 #	tst%c	%s
#	%s	 #	tst%c	%s
#	%s	 L%d
 #	incl	locprof+%d
 #L%d:
 #	incl	locprof+%d
 #	tst%c	%s
 #	jbr	L%d
 %s+%d %s %d ) #	mov%c	%s,%s
 #	pushl	%s
 #	movd	%s,%s
 #	cvt%cl	%s,%s
 #	clr%c	%s
 #	mov%c	%s,%s
 add #	.long	%s
 #	mov%c	%s,%s
 #	ashl	%s,%s,%s
 #	mov%c	%s,%s
 #	movl	%s,%s
 #	addl3	%s,%s,%s
 #	addl2	%s,%s
 #	ashl	%s,%s,%s
 #	ashl	%s,%s,%s
 #	movl	%s,%s
 sub urem #	div%c3	%s,%s,%s
 #	mul%c2	%s,%s
 #	sub%c3	%s,%s,%s
 mul %s+%d %s %d 0 bis add %s #	movl	%s,%s
 #	extzv	$%d,$%d,%s,%s
 #	subl3	%s,$32,%s
 #	extzv	%s,%s,%s,%s
 %s *%s (%s) *%s (%s)+ #	mov%c	%s,%s
 %s[%s] #	mov%c	%s,%s
 %s(%s) #	mov%c	%s,%s
 %d(%s) -(%s) (r%d)[r%d] *%s #	mov%c	%s,%s
 (%s) #	mov%c	%s,%s
 #	movl	%s,%s
 #	movl	%s,%s
 codegen failure in struct asg codgen fail in stasg #	movc3	$%d,%s,%s
 #	subl3	$%d,r3,r0
 %d(%s) %d(%s) #	mov%c	%s,%s
 #	pushal	%s
 #	mova%c	%s,%s
 ) #	mneg%c	%s,%s
 #	insv	%s,%c%d,%c%d,%s
 #	movl	%s,%s
 #	mov%c	%s,%s
  L� O� R� U� X� [� ^� a� d� g� j� n� r� v� z� ~� �� �� lbbwwllllfd??                                      ����                                     ����                                                   out of temporary trees %d(%s) %s %s %d(%s) unk mnod in copymnod #	subl2	$%d,sp
 #	subl2	$%d,r3
 #	movc3	$%d,(r3),(sp)
 #	pushl	%s
 #	movq	%s,-(sp)
 #	subl2	$%d,sp
 #	movc3	$%d,%s,(sp)
 %s #specialreg not free
 codegen: rewriting asgop fldstar
 r0 r1 r2 r3 r4 r5 r6 r7 r8 r9 r10 r11 r12 r13 r14 r15 fp ap ,D	     
   d   �  '  �� @B ���  �� ʚ;����-2147483648    @          �                  @                             0123456789abcdeflookup(%s, %d), stwart=%d, instruct=%d
 symbol table full cannot allocate hash table cannot allocate string table   �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� _                                                                                                                                                                                                                                                               �� � 
� � � no name in exname buffer too short in exname #	line %d, file %s
 L%d:
 	jbr	L%d
 #jmp L%d
 	movab	L%d,r0
 #ret %d
 	incl	locprof+%d
 	ret
 funny alignment: %d funny alignment: %d 	.align	%d
 
 
	.byte	 , 0x%x 	.long	0x%lx
  r0 r1 r2 r3 r4 r5 r6 r7 r8 r9 r10 r11 ap fp sp pc 	.text
 	.data
 	.data
 	.data	2
 	.data	1
   ttype(0%o) rbusy( %s,   )
 big register register allocation error   h� m� r� w� |� �� �� �� �� �� � prbuf overflow unexpected op in commutes -(sp) jweird ) #	moval	%s,r0
 r0 (addrsimp) rewrite struct asg hasqnode
 unk op in copytree incomprehensible type unk mnod in sideffects expression too complicated    jeql jneq jgtr jgeq jlss jleq jgtru jgequ jlssu jlequ             (((((                  H����������������������                                                                                                                                        �	 �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                $�    �������5� 4� 4� 4� 4� 2   �X	                                                                                                                                                                                 